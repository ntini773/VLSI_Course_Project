magic
tech scmos
timestamp 1732007959
<< nwell >>
rect 2237 -1471 2261 -1431
rect 2281 -1441 2318 -1439
rect 2281 -1496 2319 -1441
rect 2325 -1496 2368 -1444
rect 77 -1548 101 -1508
rect 121 -1518 158 -1516
rect 121 -1573 159 -1518
rect 165 -1573 208 -1521
rect 2236 -1563 2260 -1523
rect 76 -1640 100 -1600
rect 927 -1678 951 -1616
rect 977 -1677 1001 -1615
rect 1027 -1677 1051 -1615
rect 1074 -1677 1098 -1615
rect -284 -1756 -248 -1716
rect -242 -1763 -218 -1723
rect 2234 -1789 2258 -1749
rect 2278 -1759 2315 -1757
rect 2278 -1814 2316 -1759
rect 2322 -1814 2365 -1762
rect 90 -1894 114 -1854
rect 134 -1864 171 -1862
rect 134 -1919 172 -1864
rect 178 -1919 221 -1867
rect 1396 -1899 1420 -1847
rect 1434 -1899 1458 -1847
rect 1478 -1899 1502 -1847
rect 1516 -1899 1540 -1847
rect 1562 -1897 1586 -1845
rect 2233 -1881 2257 -1841
rect 89 -1986 113 -1946
rect -282 -2106 -246 -2066
rect -240 -2113 -216 -2073
rect 82 -2186 106 -2146
rect 126 -2156 163 -2154
rect 126 -2211 164 -2156
rect 2236 -2158 2260 -2118
rect 2280 -2128 2317 -2126
rect 170 -2211 213 -2159
rect 2280 -2183 2318 -2128
rect 2324 -2183 2367 -2131
rect 81 -2278 105 -2238
rect 2235 -2250 2259 -2210
rect -274 -2398 -238 -2358
rect -232 -2405 -208 -2365
rect 83 -2489 107 -2449
rect 127 -2459 164 -2457
rect 127 -2514 165 -2459
rect 171 -2514 214 -2462
rect 2251 -2491 2275 -2451
rect 2295 -2461 2332 -2459
rect 2295 -2516 2333 -2461
rect 2339 -2516 2382 -2464
rect 82 -2581 106 -2541
rect 2250 -2583 2274 -2543
rect -286 -2764 -250 -2724
rect -244 -2771 -220 -2731
<< ntransistor >>
rect 2248 -1489 2250 -1479
rect 88 -1566 90 -1556
rect 2295 -1546 2297 -1526
rect 2305 -1546 2307 -1526
rect 2339 -1546 2341 -1526
rect 2349 -1546 2351 -1526
rect 2247 -1581 2249 -1571
rect 135 -1623 137 -1603
rect 145 -1623 147 -1603
rect 179 -1623 181 -1603
rect 189 -1623 191 -1603
rect 87 -1658 89 -1648
rect -273 -1799 -271 -1779
rect -262 -1799 -260 -1779
rect -231 -1781 -229 -1771
rect 2245 -1807 2247 -1797
rect 101 -1912 103 -1902
rect 148 -1969 150 -1949
rect 158 -1969 160 -1949
rect 192 -1969 194 -1949
rect 202 -1969 204 -1949
rect 874 -1958 876 -1858
rect 902 -1958 904 -1858
rect 929 -1958 931 -1858
rect 968 -1958 970 -1858
rect 996 -1958 998 -1858
rect 1023 -1958 1025 -1858
rect 1063 -1957 1065 -1857
rect 1091 -1957 1093 -1857
rect 1118 -1957 1120 -1857
rect 1154 -1957 1156 -1857
rect 2292 -1864 2294 -1844
rect 2302 -1864 2304 -1844
rect 2336 -1864 2338 -1844
rect 2346 -1864 2348 -1844
rect 2244 -1899 2246 -1889
rect 1407 -1931 1409 -1911
rect 1445 -1931 1447 -1911
rect 1489 -1931 1491 -1911
rect 1527 -1931 1529 -1911
rect 1573 -1929 1575 -1909
rect 100 -2004 102 -1994
rect -271 -2149 -269 -2129
rect -260 -2149 -258 -2129
rect -229 -2131 -227 -2121
rect 93 -2204 95 -2194
rect 2247 -2176 2249 -2166
rect 140 -2261 142 -2241
rect 150 -2261 152 -2241
rect 184 -2261 186 -2241
rect 194 -2261 196 -2241
rect 2294 -2233 2296 -2213
rect 2304 -2233 2306 -2213
rect 2338 -2233 2340 -2213
rect 2348 -2233 2350 -2213
rect 2246 -2268 2248 -2258
rect 92 -2296 94 -2286
rect -263 -2441 -261 -2421
rect -252 -2441 -250 -2421
rect -221 -2423 -219 -2413
rect 94 -2507 96 -2497
rect 2262 -2509 2264 -2499
rect 141 -2564 143 -2544
rect 151 -2564 153 -2544
rect 185 -2564 187 -2544
rect 195 -2564 197 -2544
rect 2309 -2566 2311 -2546
rect 2319 -2566 2321 -2546
rect 2353 -2566 2355 -2546
rect 2363 -2566 2365 -2546
rect 93 -2599 95 -2589
rect 2261 -2601 2263 -2591
rect -275 -2807 -273 -2787
rect -264 -2807 -262 -2787
rect -233 -2789 -231 -2779
<< ptransistor >>
rect 2248 -1465 2250 -1445
rect 2295 -1490 2297 -1450
rect 2305 -1490 2307 -1450
rect 2339 -1490 2341 -1450
rect 2349 -1490 2351 -1450
rect 88 -1542 90 -1522
rect 135 -1567 137 -1527
rect 145 -1567 147 -1527
rect 179 -1567 181 -1527
rect 189 -1567 191 -1527
rect 2247 -1557 2249 -1537
rect 87 -1634 89 -1614
rect 938 -1672 940 -1622
rect 988 -1671 990 -1621
rect 1038 -1671 1040 -1621
rect 1085 -1671 1087 -1621
rect -273 -1750 -271 -1730
rect -262 -1750 -260 -1730
rect -231 -1757 -229 -1737
rect 2245 -1783 2247 -1763
rect 2292 -1808 2294 -1768
rect 2302 -1808 2304 -1768
rect 2336 -1808 2338 -1768
rect 2346 -1808 2348 -1768
rect 101 -1888 103 -1868
rect 148 -1913 150 -1873
rect 158 -1913 160 -1873
rect 192 -1913 194 -1873
rect 202 -1913 204 -1873
rect 100 -1980 102 -1960
rect 1407 -1893 1409 -1853
rect 1445 -1893 1447 -1853
rect 1489 -1893 1491 -1853
rect 1527 -1893 1529 -1853
rect 1573 -1891 1575 -1851
rect 2244 -1875 2246 -1855
rect -271 -2100 -269 -2080
rect -260 -2100 -258 -2080
rect -229 -2107 -227 -2087
rect 2247 -2152 2249 -2132
rect 93 -2180 95 -2160
rect 140 -2205 142 -2165
rect 150 -2205 152 -2165
rect 184 -2205 186 -2165
rect 194 -2205 196 -2165
rect 2294 -2177 2296 -2137
rect 2304 -2177 2306 -2137
rect 2338 -2177 2340 -2137
rect 2348 -2177 2350 -2137
rect 92 -2272 94 -2252
rect 2246 -2244 2248 -2224
rect -263 -2392 -261 -2372
rect -252 -2392 -250 -2372
rect -221 -2399 -219 -2379
rect 94 -2483 96 -2463
rect 141 -2508 143 -2468
rect 151 -2508 153 -2468
rect 185 -2508 187 -2468
rect 195 -2508 197 -2468
rect 2262 -2485 2264 -2465
rect 2309 -2510 2311 -2470
rect 2319 -2510 2321 -2470
rect 2353 -2510 2355 -2470
rect 2363 -2510 2365 -2470
rect 93 -2575 95 -2555
rect 2261 -2577 2263 -2557
rect -275 -2758 -273 -2738
rect -264 -2758 -262 -2738
rect -233 -2765 -231 -2745
<< ndiffusion >>
rect 2247 -1489 2248 -1479
rect 2250 -1489 2251 -1479
rect 87 -1566 88 -1556
rect 90 -1566 91 -1556
rect 2294 -1546 2295 -1526
rect 2297 -1546 2305 -1526
rect 2307 -1546 2308 -1526
rect 2338 -1546 2339 -1526
rect 2341 -1546 2349 -1526
rect 2351 -1546 2352 -1526
rect 2246 -1581 2247 -1571
rect 2249 -1581 2250 -1571
rect 134 -1623 135 -1603
rect 137 -1623 145 -1603
rect 147 -1623 148 -1603
rect 178 -1623 179 -1603
rect 181 -1623 189 -1603
rect 191 -1623 192 -1603
rect 86 -1658 87 -1648
rect 89 -1658 90 -1648
rect -274 -1799 -273 -1779
rect -271 -1799 -262 -1779
rect -260 -1799 -259 -1779
rect -232 -1781 -231 -1771
rect -229 -1781 -228 -1771
rect 2244 -1807 2245 -1797
rect 2247 -1807 2248 -1797
rect 100 -1912 101 -1902
rect 103 -1912 104 -1902
rect 147 -1969 148 -1949
rect 150 -1969 158 -1949
rect 160 -1969 161 -1949
rect 191 -1969 192 -1949
rect 194 -1969 202 -1949
rect 204 -1969 205 -1949
rect 873 -1958 874 -1858
rect 876 -1958 877 -1858
rect 901 -1958 902 -1858
rect 904 -1958 905 -1858
rect 928 -1958 929 -1858
rect 931 -1958 932 -1858
rect 967 -1958 968 -1858
rect 970 -1958 971 -1858
rect 995 -1958 996 -1858
rect 998 -1958 999 -1858
rect 1022 -1958 1023 -1858
rect 1025 -1958 1026 -1858
rect 1062 -1957 1063 -1857
rect 1065 -1957 1066 -1857
rect 1090 -1957 1091 -1857
rect 1093 -1957 1094 -1857
rect 1117 -1957 1118 -1857
rect 1120 -1957 1121 -1857
rect 1153 -1957 1154 -1857
rect 1156 -1957 1157 -1857
rect 2291 -1864 2292 -1844
rect 2294 -1864 2302 -1844
rect 2304 -1864 2305 -1844
rect 2335 -1864 2336 -1844
rect 2338 -1864 2346 -1844
rect 2348 -1864 2349 -1844
rect 2243 -1899 2244 -1889
rect 2246 -1899 2247 -1889
rect 1406 -1931 1407 -1911
rect 1409 -1931 1410 -1911
rect 1444 -1931 1445 -1911
rect 1447 -1931 1448 -1911
rect 1488 -1931 1489 -1911
rect 1491 -1931 1492 -1911
rect 1526 -1931 1527 -1911
rect 1529 -1931 1530 -1911
rect 1572 -1929 1573 -1909
rect 1575 -1929 1576 -1909
rect 99 -2004 100 -1994
rect 102 -2004 103 -1994
rect -272 -2149 -271 -2129
rect -269 -2149 -260 -2129
rect -258 -2149 -257 -2129
rect -230 -2131 -229 -2121
rect -227 -2131 -226 -2121
rect 92 -2204 93 -2194
rect 95 -2204 96 -2194
rect 2246 -2176 2247 -2166
rect 2249 -2176 2250 -2166
rect 139 -2261 140 -2241
rect 142 -2261 150 -2241
rect 152 -2261 153 -2241
rect 183 -2261 184 -2241
rect 186 -2261 194 -2241
rect 196 -2261 197 -2241
rect 2293 -2233 2294 -2213
rect 2296 -2233 2304 -2213
rect 2306 -2233 2307 -2213
rect 2337 -2233 2338 -2213
rect 2340 -2233 2348 -2213
rect 2350 -2233 2351 -2213
rect 2245 -2268 2246 -2258
rect 2248 -2268 2249 -2258
rect 91 -2296 92 -2286
rect 94 -2296 95 -2286
rect -264 -2441 -263 -2421
rect -261 -2441 -252 -2421
rect -250 -2441 -249 -2421
rect -222 -2423 -221 -2413
rect -219 -2423 -218 -2413
rect 93 -2507 94 -2497
rect 96 -2507 97 -2497
rect 2261 -2509 2262 -2499
rect 2264 -2509 2265 -2499
rect 140 -2564 141 -2544
rect 143 -2564 151 -2544
rect 153 -2564 154 -2544
rect 184 -2564 185 -2544
rect 187 -2564 195 -2544
rect 197 -2564 198 -2544
rect 2308 -2566 2309 -2546
rect 2311 -2566 2319 -2546
rect 2321 -2566 2322 -2546
rect 2352 -2566 2353 -2546
rect 2355 -2566 2363 -2546
rect 2365 -2566 2366 -2546
rect 92 -2599 93 -2589
rect 95 -2599 96 -2589
rect 2260 -2601 2261 -2591
rect 2263 -2601 2264 -2591
rect -276 -2807 -275 -2787
rect -273 -2807 -264 -2787
rect -262 -2807 -261 -2787
rect -234 -2789 -233 -2779
rect -231 -2789 -230 -2779
<< pdiffusion >>
rect 2247 -1465 2248 -1445
rect 2250 -1465 2251 -1445
rect 2294 -1490 2295 -1450
rect 2297 -1490 2299 -1450
rect 2303 -1490 2305 -1450
rect 2307 -1490 2308 -1450
rect 2338 -1490 2339 -1450
rect 2341 -1490 2343 -1450
rect 2347 -1490 2349 -1450
rect 2351 -1490 2352 -1450
rect 87 -1542 88 -1522
rect 90 -1542 91 -1522
rect 134 -1567 135 -1527
rect 137 -1567 139 -1527
rect 143 -1567 145 -1527
rect 147 -1567 148 -1527
rect 178 -1567 179 -1527
rect 181 -1567 183 -1527
rect 187 -1567 189 -1527
rect 191 -1567 192 -1527
rect 2246 -1557 2247 -1537
rect 2249 -1557 2250 -1537
rect 86 -1634 87 -1614
rect 89 -1634 90 -1614
rect 937 -1672 938 -1622
rect 940 -1672 941 -1622
rect 987 -1671 988 -1621
rect 990 -1671 991 -1621
rect 1037 -1671 1038 -1621
rect 1040 -1671 1041 -1621
rect 1084 -1671 1085 -1621
rect 1087 -1671 1088 -1621
rect -274 -1750 -273 -1730
rect -271 -1750 -267 -1730
rect -263 -1750 -262 -1730
rect -260 -1750 -259 -1730
rect -232 -1757 -231 -1737
rect -229 -1757 -228 -1737
rect 2244 -1783 2245 -1763
rect 2247 -1783 2248 -1763
rect 2291 -1808 2292 -1768
rect 2294 -1808 2296 -1768
rect 2300 -1808 2302 -1768
rect 2304 -1808 2305 -1768
rect 2335 -1808 2336 -1768
rect 2338 -1808 2340 -1768
rect 2344 -1808 2346 -1768
rect 2348 -1808 2349 -1768
rect 100 -1888 101 -1868
rect 103 -1888 104 -1868
rect 147 -1913 148 -1873
rect 150 -1913 152 -1873
rect 156 -1913 158 -1873
rect 160 -1913 161 -1873
rect 191 -1913 192 -1873
rect 194 -1913 196 -1873
rect 200 -1913 202 -1873
rect 204 -1913 205 -1873
rect 99 -1980 100 -1960
rect 102 -1980 103 -1960
rect 1406 -1893 1407 -1853
rect 1409 -1893 1410 -1853
rect 1444 -1893 1445 -1853
rect 1447 -1893 1448 -1853
rect 1488 -1893 1489 -1853
rect 1491 -1893 1492 -1853
rect 1526 -1893 1527 -1853
rect 1529 -1893 1530 -1853
rect 1572 -1891 1573 -1851
rect 1575 -1891 1576 -1851
rect 2243 -1875 2244 -1855
rect 2246 -1875 2247 -1855
rect -272 -2100 -271 -2080
rect -269 -2100 -265 -2080
rect -261 -2100 -260 -2080
rect -258 -2100 -257 -2080
rect -230 -2107 -229 -2087
rect -227 -2107 -226 -2087
rect 2246 -2152 2247 -2132
rect 2249 -2152 2250 -2132
rect 92 -2180 93 -2160
rect 95 -2180 96 -2160
rect 139 -2205 140 -2165
rect 142 -2205 144 -2165
rect 148 -2205 150 -2165
rect 152 -2205 153 -2165
rect 183 -2205 184 -2165
rect 186 -2205 188 -2165
rect 192 -2205 194 -2165
rect 196 -2205 197 -2165
rect 2293 -2177 2294 -2137
rect 2296 -2177 2298 -2137
rect 2302 -2177 2304 -2137
rect 2306 -2177 2307 -2137
rect 2337 -2177 2338 -2137
rect 2340 -2177 2342 -2137
rect 2346 -2177 2348 -2137
rect 2350 -2177 2351 -2137
rect 91 -2272 92 -2252
rect 94 -2272 95 -2252
rect 2245 -2244 2246 -2224
rect 2248 -2244 2249 -2224
rect -264 -2392 -263 -2372
rect -261 -2392 -257 -2372
rect -253 -2392 -252 -2372
rect -250 -2392 -249 -2372
rect -222 -2399 -221 -2379
rect -219 -2399 -218 -2379
rect 93 -2483 94 -2463
rect 96 -2483 97 -2463
rect 140 -2508 141 -2468
rect 143 -2508 145 -2468
rect 149 -2508 151 -2468
rect 153 -2508 154 -2468
rect 184 -2508 185 -2468
rect 187 -2508 189 -2468
rect 193 -2508 195 -2468
rect 197 -2508 198 -2468
rect 2261 -2485 2262 -2465
rect 2264 -2485 2265 -2465
rect 2308 -2510 2309 -2470
rect 2311 -2510 2313 -2470
rect 2317 -2510 2319 -2470
rect 2321 -2510 2322 -2470
rect 2352 -2510 2353 -2470
rect 2355 -2510 2357 -2470
rect 2361 -2510 2363 -2470
rect 2365 -2510 2366 -2470
rect 92 -2575 93 -2555
rect 95 -2575 96 -2555
rect 2260 -2577 2261 -2557
rect 2263 -2577 2264 -2557
rect -276 -2758 -275 -2738
rect -273 -2758 -269 -2738
rect -265 -2758 -264 -2738
rect -262 -2758 -261 -2738
rect -234 -2765 -233 -2745
rect -231 -2765 -230 -2745
<< ndcontact >>
rect 2243 -1489 2247 -1479
rect 2251 -1489 2255 -1479
rect 83 -1566 87 -1556
rect 91 -1566 95 -1556
rect 2290 -1546 2294 -1526
rect 2308 -1546 2312 -1526
rect 2334 -1546 2338 -1526
rect 2352 -1546 2356 -1526
rect 2242 -1581 2246 -1571
rect 2250 -1581 2254 -1571
rect 130 -1623 134 -1603
rect 148 -1623 152 -1603
rect 174 -1623 178 -1603
rect 192 -1623 196 -1603
rect 82 -1658 86 -1648
rect 90 -1658 94 -1648
rect -278 -1799 -274 -1779
rect -259 -1799 -255 -1779
rect -236 -1781 -232 -1771
rect -228 -1781 -224 -1771
rect 2240 -1807 2244 -1797
rect 2248 -1807 2252 -1797
rect 96 -1912 100 -1902
rect 104 -1912 108 -1902
rect 143 -1969 147 -1949
rect 161 -1969 165 -1949
rect 187 -1969 191 -1949
rect 205 -1969 209 -1949
rect 869 -1958 873 -1858
rect 877 -1958 881 -1858
rect 897 -1958 901 -1858
rect 905 -1958 909 -1858
rect 924 -1958 928 -1858
rect 932 -1958 936 -1858
rect 963 -1958 967 -1858
rect 971 -1958 975 -1858
rect 991 -1958 995 -1858
rect 999 -1958 1003 -1858
rect 1018 -1958 1022 -1858
rect 1026 -1958 1030 -1858
rect 1058 -1957 1062 -1857
rect 1066 -1957 1070 -1857
rect 1086 -1957 1090 -1857
rect 1094 -1957 1098 -1857
rect 1113 -1957 1117 -1857
rect 1121 -1957 1125 -1857
rect 1149 -1957 1153 -1857
rect 1157 -1957 1161 -1857
rect 2287 -1864 2291 -1844
rect 2305 -1864 2309 -1844
rect 2331 -1864 2335 -1844
rect 2349 -1864 2353 -1844
rect 2239 -1899 2243 -1889
rect 2247 -1899 2251 -1889
rect 1402 -1931 1406 -1911
rect 1410 -1931 1414 -1911
rect 1440 -1931 1444 -1911
rect 1448 -1931 1452 -1911
rect 1484 -1931 1488 -1911
rect 1492 -1931 1496 -1911
rect 1522 -1931 1526 -1911
rect 1530 -1931 1534 -1911
rect 1568 -1929 1572 -1909
rect 1576 -1929 1580 -1909
rect 95 -2004 99 -1994
rect 103 -2004 107 -1994
rect -276 -2149 -272 -2129
rect -257 -2149 -253 -2129
rect -234 -2131 -230 -2121
rect -226 -2131 -222 -2121
rect 88 -2204 92 -2194
rect 96 -2204 100 -2194
rect 2242 -2176 2246 -2166
rect 2250 -2176 2254 -2166
rect 135 -2261 139 -2241
rect 153 -2261 157 -2241
rect 179 -2261 183 -2241
rect 197 -2261 201 -2241
rect 2289 -2233 2293 -2213
rect 2307 -2233 2311 -2213
rect 2333 -2233 2337 -2213
rect 2351 -2233 2355 -2213
rect 2241 -2268 2245 -2258
rect 2249 -2268 2253 -2258
rect 87 -2296 91 -2286
rect 95 -2296 99 -2286
rect -268 -2441 -264 -2421
rect -249 -2441 -245 -2421
rect -226 -2423 -222 -2413
rect -218 -2423 -214 -2413
rect 89 -2507 93 -2497
rect 97 -2507 101 -2497
rect 2257 -2509 2261 -2499
rect 2265 -2509 2269 -2499
rect 136 -2564 140 -2544
rect 154 -2564 158 -2544
rect 180 -2564 184 -2544
rect 198 -2564 202 -2544
rect 2304 -2566 2308 -2546
rect 2322 -2566 2326 -2546
rect 2348 -2566 2352 -2546
rect 2366 -2566 2370 -2546
rect 88 -2599 92 -2589
rect 96 -2599 100 -2589
rect 2256 -2601 2260 -2591
rect 2264 -2601 2268 -2591
rect -280 -2807 -276 -2787
rect -261 -2807 -257 -2787
rect -238 -2789 -234 -2779
rect -230 -2789 -226 -2779
<< pdcontact >>
rect 2243 -1465 2247 -1445
rect 2251 -1465 2255 -1445
rect 2290 -1490 2294 -1450
rect 2299 -1490 2303 -1450
rect 2308 -1490 2312 -1450
rect 2334 -1490 2338 -1450
rect 2343 -1490 2347 -1450
rect 2352 -1490 2356 -1450
rect 83 -1542 87 -1522
rect 91 -1542 95 -1522
rect 130 -1567 134 -1527
rect 139 -1567 143 -1527
rect 148 -1567 152 -1527
rect 174 -1567 178 -1527
rect 183 -1567 187 -1527
rect 192 -1567 196 -1527
rect 2242 -1557 2246 -1537
rect 2250 -1557 2254 -1537
rect 82 -1634 86 -1614
rect 90 -1634 94 -1614
rect 933 -1672 937 -1622
rect 941 -1672 945 -1622
rect 983 -1671 987 -1621
rect 991 -1671 995 -1621
rect 1033 -1671 1037 -1621
rect 1041 -1671 1045 -1621
rect 1080 -1671 1084 -1621
rect 1088 -1671 1092 -1621
rect -278 -1750 -274 -1730
rect -267 -1750 -263 -1730
rect -259 -1750 -255 -1730
rect -236 -1757 -232 -1737
rect -228 -1757 -224 -1737
rect 2240 -1783 2244 -1763
rect 2248 -1783 2252 -1763
rect 2287 -1808 2291 -1768
rect 2296 -1808 2300 -1768
rect 2305 -1808 2309 -1768
rect 2331 -1808 2335 -1768
rect 2340 -1808 2344 -1768
rect 2349 -1808 2353 -1768
rect 96 -1888 100 -1868
rect 104 -1888 108 -1868
rect 143 -1913 147 -1873
rect 152 -1913 156 -1873
rect 161 -1913 165 -1873
rect 187 -1913 191 -1873
rect 196 -1913 200 -1873
rect 205 -1913 209 -1873
rect 95 -1980 99 -1960
rect 103 -1980 107 -1960
rect 1402 -1893 1406 -1853
rect 1410 -1893 1414 -1853
rect 1440 -1893 1444 -1853
rect 1448 -1893 1452 -1853
rect 1484 -1893 1488 -1853
rect 1492 -1893 1496 -1853
rect 1522 -1893 1526 -1853
rect 1530 -1893 1534 -1853
rect 1568 -1891 1572 -1851
rect 1576 -1891 1580 -1851
rect 2239 -1875 2243 -1855
rect 2247 -1875 2251 -1855
rect -276 -2100 -272 -2080
rect -265 -2100 -261 -2080
rect -257 -2100 -253 -2080
rect -234 -2107 -230 -2087
rect -226 -2107 -222 -2087
rect 2242 -2152 2246 -2132
rect 2250 -2152 2254 -2132
rect 88 -2180 92 -2160
rect 96 -2180 100 -2160
rect 135 -2205 139 -2165
rect 144 -2205 148 -2165
rect 153 -2205 157 -2165
rect 179 -2205 183 -2165
rect 188 -2205 192 -2165
rect 197 -2205 201 -2165
rect 2289 -2177 2293 -2137
rect 2298 -2177 2302 -2137
rect 2307 -2177 2311 -2137
rect 2333 -2177 2337 -2137
rect 2342 -2177 2346 -2137
rect 2351 -2177 2355 -2137
rect 87 -2272 91 -2252
rect 95 -2272 99 -2252
rect 2241 -2244 2245 -2224
rect 2249 -2244 2253 -2224
rect -268 -2392 -264 -2372
rect -257 -2392 -253 -2372
rect -249 -2392 -245 -2372
rect -226 -2399 -222 -2379
rect -218 -2399 -214 -2379
rect 89 -2483 93 -2463
rect 97 -2483 101 -2463
rect 136 -2508 140 -2468
rect 145 -2508 149 -2468
rect 154 -2508 158 -2468
rect 180 -2508 184 -2468
rect 189 -2508 193 -2468
rect 198 -2508 202 -2468
rect 2257 -2485 2261 -2465
rect 2265 -2485 2269 -2465
rect 2304 -2510 2308 -2470
rect 2313 -2510 2317 -2470
rect 2322 -2510 2326 -2470
rect 2348 -2510 2352 -2470
rect 2357 -2510 2361 -2470
rect 2366 -2510 2370 -2470
rect 88 -2575 92 -2555
rect 96 -2575 100 -2555
rect 2256 -2577 2260 -2557
rect 2264 -2577 2268 -2557
rect -280 -2758 -276 -2738
rect -269 -2758 -265 -2738
rect -261 -2758 -257 -2738
rect -238 -2765 -234 -2745
rect -230 -2765 -226 -2745
<< psubstratepcontact >>
rect 2257 -1498 2262 -1494
rect 2322 -1553 2330 -1549
rect 97 -1575 102 -1571
rect 2256 -1590 2261 -1586
rect 162 -1630 170 -1626
rect 96 -1667 101 -1663
rect -222 -1790 -217 -1786
rect 2254 -1816 2259 -1812
rect 110 -1921 115 -1917
rect 2319 -1871 2327 -1867
rect 2253 -1908 2258 -1904
rect 175 -1976 183 -1972
rect 109 -2013 114 -2009
rect -220 -2140 -215 -2136
rect 2256 -2185 2261 -2181
rect 102 -2213 107 -2209
rect 2321 -2240 2329 -2236
rect 167 -2268 175 -2264
rect 2255 -2277 2260 -2273
rect 101 -2305 106 -2301
rect -212 -2432 -207 -2428
rect 103 -2516 108 -2512
rect 2271 -2518 2276 -2514
rect 168 -2571 176 -2567
rect 2336 -2573 2344 -2569
rect 102 -2608 107 -2604
rect 2270 -2610 2275 -2606
rect -224 -2798 -219 -2794
<< nsubstratencontact >>
rect 2253 -1438 2257 -1434
rect 2289 -1446 2295 -1442
rect 2360 -1452 2365 -1447
rect 93 -1515 97 -1511
rect 129 -1523 135 -1519
rect 200 -1529 205 -1524
rect 2252 -1530 2256 -1526
rect 92 -1607 96 -1603
rect 928 -1616 932 -1611
rect 978 -1615 982 -1610
rect 1028 -1615 1032 -1610
rect 1075 -1615 1079 -1610
rect -278 -1725 -274 -1719
rect -226 -1730 -222 -1726
rect 2250 -1756 2254 -1752
rect 2286 -1764 2292 -1760
rect 2357 -1770 2362 -1765
rect 1397 -1847 1401 -1843
rect 1435 -1847 1439 -1843
rect 1479 -1847 1483 -1843
rect 1517 -1847 1521 -1843
rect 1563 -1845 1567 -1841
rect 2249 -1848 2253 -1844
rect 106 -1861 110 -1857
rect 142 -1869 148 -1865
rect 213 -1875 218 -1870
rect 105 -1953 109 -1949
rect -276 -2075 -272 -2069
rect -224 -2080 -220 -2076
rect 2252 -2125 2256 -2121
rect 98 -2153 102 -2149
rect 2288 -2133 2294 -2129
rect 134 -2161 140 -2157
rect 205 -2167 210 -2162
rect 2359 -2139 2364 -2134
rect 2251 -2217 2255 -2213
rect 97 -2245 101 -2241
rect -268 -2367 -264 -2361
rect -216 -2372 -212 -2368
rect 99 -2456 103 -2452
rect 2267 -2458 2271 -2454
rect 135 -2464 141 -2460
rect 206 -2470 211 -2465
rect 2303 -2466 2309 -2462
rect 2374 -2472 2379 -2467
rect 98 -2548 102 -2544
rect 2266 -2550 2270 -2546
rect -280 -2733 -276 -2727
rect -228 -2738 -224 -2734
<< polysilicon >>
rect 2248 -1445 2250 -1441
rect 2295 -1450 2297 -1447
rect 2305 -1450 2307 -1447
rect 2339 -1450 2341 -1447
rect 2349 -1450 2351 -1447
rect 2248 -1479 2250 -1465
rect 2248 -1492 2250 -1489
rect 2295 -1494 2297 -1490
rect 2296 -1499 2297 -1494
rect 88 -1522 90 -1518
rect 135 -1527 137 -1524
rect 145 -1527 147 -1524
rect 179 -1527 181 -1524
rect 189 -1527 191 -1524
rect 88 -1556 90 -1542
rect 88 -1569 90 -1566
rect 2295 -1526 2297 -1499
rect 2305 -1518 2307 -1490
rect 2305 -1526 2307 -1522
rect 2339 -1526 2341 -1490
rect 2349 -1526 2351 -1490
rect 2247 -1537 2249 -1533
rect 2295 -1549 2297 -1546
rect 2305 -1549 2307 -1546
rect 2339 -1549 2341 -1546
rect 2349 -1549 2351 -1546
rect 135 -1571 137 -1567
rect 136 -1576 137 -1571
rect 135 -1603 137 -1576
rect 145 -1595 147 -1567
rect 145 -1603 147 -1599
rect 179 -1603 181 -1567
rect 189 -1603 191 -1567
rect 2247 -1571 2249 -1557
rect 2247 -1584 2249 -1581
rect 87 -1614 89 -1610
rect 938 -1622 940 -1619
rect 988 -1621 990 -1618
rect 1038 -1621 1040 -1618
rect 1085 -1621 1087 -1618
rect 135 -1626 137 -1623
rect 145 -1626 147 -1623
rect 179 -1626 181 -1623
rect 189 -1626 191 -1623
rect 87 -1648 89 -1634
rect 87 -1661 89 -1658
rect 938 -1695 940 -1672
rect 988 -1694 990 -1671
rect 1038 -1694 1040 -1671
rect 1085 -1694 1087 -1671
rect -273 -1730 -271 -1727
rect -262 -1730 -260 -1727
rect -231 -1737 -229 -1733
rect -273 -1779 -271 -1750
rect -262 -1779 -260 -1750
rect -231 -1771 -229 -1757
rect 2245 -1763 2247 -1759
rect -231 -1784 -229 -1781
rect 2292 -1768 2294 -1765
rect 2302 -1768 2304 -1765
rect 2336 -1768 2338 -1765
rect 2346 -1768 2348 -1765
rect 2245 -1797 2247 -1783
rect -273 -1802 -271 -1799
rect -262 -1802 -260 -1799
rect 2245 -1810 2247 -1807
rect 2292 -1812 2294 -1808
rect 2293 -1817 2294 -1812
rect 2292 -1844 2294 -1817
rect 2302 -1836 2304 -1808
rect 2302 -1844 2304 -1840
rect 2336 -1844 2338 -1808
rect 2346 -1844 2348 -1808
rect 1407 -1853 1409 -1850
rect 1445 -1853 1447 -1850
rect 1489 -1853 1491 -1850
rect 1527 -1853 1529 -1850
rect 1573 -1851 1575 -1848
rect 874 -1858 876 -1855
rect 902 -1858 904 -1855
rect 929 -1858 931 -1855
rect 968 -1858 970 -1855
rect 996 -1858 998 -1855
rect 1023 -1858 1025 -1855
rect 1063 -1857 1065 -1854
rect 1091 -1857 1093 -1854
rect 1118 -1857 1120 -1854
rect 1154 -1857 1156 -1854
rect 101 -1868 103 -1864
rect 148 -1873 150 -1870
rect 158 -1873 160 -1870
rect 192 -1873 194 -1870
rect 202 -1873 204 -1870
rect 101 -1902 103 -1888
rect 101 -1915 103 -1912
rect 148 -1917 150 -1913
rect 149 -1922 150 -1917
rect 148 -1949 150 -1922
rect 158 -1941 160 -1913
rect 158 -1949 160 -1945
rect 192 -1949 194 -1913
rect 202 -1949 204 -1913
rect 100 -1960 102 -1956
rect 2244 -1855 2246 -1851
rect 2292 -1867 2294 -1864
rect 2302 -1867 2304 -1864
rect 2336 -1867 2338 -1864
rect 2346 -1867 2348 -1864
rect 2244 -1889 2246 -1875
rect 1407 -1911 1409 -1893
rect 1445 -1911 1447 -1893
rect 1489 -1911 1491 -1893
rect 1527 -1911 1529 -1893
rect 1573 -1909 1575 -1891
rect 2244 -1902 2246 -1899
rect 1407 -1935 1409 -1931
rect 1445 -1935 1447 -1931
rect 1489 -1935 1491 -1931
rect 1527 -1935 1529 -1931
rect 1573 -1933 1575 -1929
rect 148 -1972 150 -1969
rect 158 -1972 160 -1969
rect 192 -1972 194 -1969
rect 202 -1972 204 -1969
rect 874 -1970 876 -1958
rect 902 -1970 904 -1958
rect 929 -1970 931 -1958
rect 968 -1970 970 -1958
rect 996 -1970 998 -1958
rect 1023 -1970 1025 -1958
rect 1063 -1969 1065 -1957
rect 1091 -1969 1093 -1957
rect 1118 -1969 1120 -1957
rect 1154 -1969 1156 -1957
rect 100 -1994 102 -1980
rect 100 -2007 102 -2004
rect -271 -2080 -269 -2077
rect -260 -2080 -258 -2077
rect -229 -2087 -227 -2083
rect -271 -2129 -269 -2100
rect -260 -2129 -258 -2100
rect -229 -2121 -227 -2107
rect -229 -2134 -227 -2131
rect 2247 -2132 2249 -2128
rect -271 -2152 -269 -2149
rect -260 -2152 -258 -2149
rect 2294 -2137 2296 -2134
rect 2304 -2137 2306 -2134
rect 2338 -2137 2340 -2134
rect 2348 -2137 2350 -2134
rect 93 -2160 95 -2156
rect 140 -2165 142 -2162
rect 150 -2165 152 -2162
rect 184 -2165 186 -2162
rect 194 -2165 196 -2162
rect 93 -2194 95 -2180
rect 93 -2207 95 -2204
rect 2247 -2166 2249 -2152
rect 2247 -2179 2249 -2176
rect 2294 -2181 2296 -2177
rect 2295 -2186 2296 -2181
rect 140 -2209 142 -2205
rect 141 -2214 142 -2209
rect 140 -2241 142 -2214
rect 150 -2233 152 -2205
rect 150 -2241 152 -2237
rect 184 -2241 186 -2205
rect 194 -2241 196 -2205
rect 2294 -2213 2296 -2186
rect 2304 -2205 2306 -2177
rect 2304 -2213 2306 -2209
rect 2338 -2213 2340 -2177
rect 2348 -2213 2350 -2177
rect 2246 -2224 2248 -2220
rect 92 -2252 94 -2248
rect 2294 -2236 2296 -2233
rect 2304 -2236 2306 -2233
rect 2338 -2236 2340 -2233
rect 2348 -2236 2350 -2233
rect 2246 -2258 2248 -2244
rect 140 -2264 142 -2261
rect 150 -2264 152 -2261
rect 184 -2264 186 -2261
rect 194 -2264 196 -2261
rect 2246 -2271 2248 -2268
rect 92 -2286 94 -2272
rect 92 -2299 94 -2296
rect -263 -2372 -261 -2369
rect -252 -2372 -250 -2369
rect -221 -2379 -219 -2375
rect -263 -2421 -261 -2392
rect -252 -2421 -250 -2392
rect -221 -2413 -219 -2399
rect -221 -2426 -219 -2423
rect -263 -2444 -261 -2441
rect -252 -2444 -250 -2441
rect 94 -2463 96 -2459
rect 2262 -2465 2264 -2461
rect 141 -2468 143 -2465
rect 151 -2468 153 -2465
rect 185 -2468 187 -2465
rect 195 -2468 197 -2465
rect 94 -2497 96 -2483
rect 94 -2510 96 -2507
rect 2309 -2470 2311 -2467
rect 2319 -2470 2321 -2467
rect 2353 -2470 2355 -2467
rect 2363 -2470 2365 -2467
rect 2262 -2499 2264 -2485
rect 141 -2512 143 -2508
rect 142 -2517 143 -2512
rect 141 -2544 143 -2517
rect 151 -2536 153 -2508
rect 151 -2544 153 -2540
rect 185 -2544 187 -2508
rect 195 -2544 197 -2508
rect 2262 -2512 2264 -2509
rect 2309 -2514 2311 -2510
rect 2310 -2519 2311 -2514
rect 93 -2555 95 -2551
rect 2309 -2546 2311 -2519
rect 2319 -2538 2321 -2510
rect 2319 -2546 2321 -2542
rect 2353 -2546 2355 -2510
rect 2363 -2546 2365 -2510
rect 2261 -2557 2263 -2553
rect 141 -2567 143 -2564
rect 151 -2567 153 -2564
rect 185 -2567 187 -2564
rect 195 -2567 197 -2564
rect 93 -2589 95 -2575
rect 2309 -2569 2311 -2566
rect 2319 -2569 2321 -2566
rect 2353 -2569 2355 -2566
rect 2363 -2569 2365 -2566
rect 2261 -2591 2263 -2577
rect 93 -2602 95 -2599
rect 2261 -2604 2263 -2601
rect -275 -2738 -273 -2735
rect -264 -2738 -262 -2735
rect -233 -2745 -231 -2741
rect -275 -2787 -273 -2758
rect -264 -2787 -262 -2758
rect -233 -2779 -231 -2765
rect -233 -2792 -231 -2789
rect -275 -2810 -273 -2807
rect -264 -2810 -262 -2807
<< polycontact >>
rect 2244 -1476 2248 -1472
rect 84 -1553 88 -1549
rect 2335 -1507 2339 -1503
rect 2345 -1515 2349 -1511
rect 175 -1584 179 -1580
rect 185 -1592 189 -1588
rect 2243 -1568 2247 -1564
rect 83 -1645 87 -1641
rect -277 -1776 -273 -1772
rect -266 -1769 -262 -1765
rect -235 -1768 -231 -1764
rect 2241 -1794 2245 -1790
rect 2332 -1825 2336 -1821
rect 2342 -1833 2346 -1829
rect 97 -1899 101 -1895
rect 188 -1930 192 -1926
rect 198 -1938 202 -1934
rect 2240 -1886 2244 -1882
rect 96 -1991 100 -1987
rect -275 -2126 -271 -2122
rect -264 -2119 -260 -2115
rect -233 -2118 -229 -2114
rect 89 -2191 93 -2187
rect 2243 -2163 2247 -2159
rect 180 -2222 184 -2218
rect 190 -2230 194 -2226
rect 2334 -2194 2338 -2190
rect 2344 -2202 2348 -2198
rect 2242 -2255 2246 -2251
rect 88 -2283 92 -2279
rect -267 -2418 -263 -2414
rect -256 -2411 -252 -2407
rect -225 -2410 -221 -2406
rect 90 -2494 94 -2490
rect 2258 -2496 2262 -2492
rect 181 -2525 185 -2521
rect 191 -2533 195 -2529
rect 2349 -2527 2353 -2523
rect 2359 -2535 2363 -2531
rect 89 -2586 93 -2582
rect 2257 -2588 2261 -2584
rect -279 -2784 -275 -2780
rect -268 -2777 -264 -2773
rect -237 -2776 -233 -2772
<< metal1 >>
rect 2241 -1434 2280 -1433
rect 2241 -1438 2253 -1434
rect 2257 -1438 2363 -1434
rect 2241 -1440 2261 -1438
rect 2243 -1445 2247 -1440
rect 2289 -1442 2294 -1438
rect 2289 -1448 2294 -1446
rect 2251 -1472 2255 -1465
rect 2290 -1450 2294 -1448
rect 2308 -1450 2312 -1438
rect 2235 -1476 2244 -1472
rect 2251 -1476 2272 -1472
rect 2251 -1479 2255 -1476
rect 2243 -1493 2247 -1489
rect 2237 -1494 2262 -1493
rect 2237 -1496 2257 -1494
rect 2237 -1499 2250 -1496
rect 2256 -1498 2257 -1496
rect 2256 -1499 2262 -1498
rect 2268 -1503 2272 -1476
rect 2334 -1444 2356 -1441
rect 2334 -1450 2338 -1444
rect 2352 -1450 2356 -1444
rect 2299 -1494 2303 -1490
rect 2334 -1494 2338 -1490
rect 2299 -1498 2338 -1494
rect 2359 -1447 2363 -1438
rect 2359 -1452 2360 -1447
rect 2343 -1496 2347 -1490
rect 2343 -1500 2360 -1496
rect 2268 -1507 2335 -1503
rect 81 -1511 120 -1510
rect 81 -1515 93 -1511
rect 97 -1515 203 -1511
rect 81 -1517 101 -1515
rect 83 -1522 87 -1517
rect 129 -1519 134 -1515
rect 129 -1525 134 -1523
rect 91 -1549 95 -1542
rect 130 -1527 134 -1525
rect 148 -1527 152 -1515
rect 75 -1553 84 -1549
rect 91 -1553 112 -1549
rect 91 -1556 95 -1553
rect 83 -1570 87 -1566
rect 77 -1571 102 -1570
rect 77 -1573 97 -1571
rect 77 -1576 90 -1573
rect 96 -1575 97 -1573
rect 96 -1576 102 -1575
rect 108 -1580 112 -1553
rect 174 -1521 196 -1518
rect 174 -1527 178 -1521
rect 192 -1527 196 -1521
rect 139 -1571 143 -1567
rect 174 -1571 178 -1567
rect 139 -1575 178 -1571
rect 199 -1524 203 -1515
rect 2272 -1515 2345 -1511
rect 199 -1529 200 -1524
rect 2241 -1526 2260 -1525
rect 2241 -1530 2252 -1526
rect 2256 -1530 2260 -1526
rect 2241 -1532 2260 -1530
rect 2242 -1537 2246 -1532
rect 183 -1573 187 -1567
rect 2250 -1564 2254 -1557
rect 2272 -1564 2276 -1515
rect 2356 -1519 2360 -1500
rect 2322 -1523 2360 -1519
rect 2322 -1526 2326 -1523
rect 2233 -1568 2243 -1564
rect 2250 -1568 2276 -1564
rect 2312 -1530 2334 -1526
rect 2290 -1549 2294 -1546
rect 2352 -1549 2356 -1546
rect 2290 -1553 2322 -1549
rect 2330 -1553 2356 -1549
rect 2250 -1571 2254 -1568
rect 183 -1577 200 -1573
rect 108 -1584 175 -1580
rect 112 -1592 185 -1588
rect 81 -1603 100 -1602
rect 81 -1607 92 -1603
rect 96 -1607 100 -1603
rect 81 -1609 100 -1607
rect 82 -1614 86 -1609
rect 90 -1641 94 -1634
rect 112 -1641 116 -1592
rect 196 -1596 200 -1577
rect 2242 -1585 2246 -1581
rect 2290 -1585 2294 -1553
rect 2236 -1586 2264 -1585
rect 2236 -1590 2256 -1586
rect 2261 -1589 2264 -1586
rect 2269 -1589 2294 -1585
rect 2236 -1591 2261 -1590
rect 162 -1600 200 -1596
rect 162 -1603 166 -1600
rect 73 -1645 83 -1641
rect 90 -1645 116 -1641
rect 152 -1607 174 -1603
rect 933 -1611 937 -1602
rect 983 -1610 987 -1601
rect 1033 -1610 1037 -1601
rect 1080 -1610 1084 -1601
rect 927 -1616 928 -1611
rect 932 -1616 951 -1611
rect 977 -1615 978 -1610
rect 982 -1615 1001 -1610
rect 1027 -1615 1028 -1610
rect 1032 -1615 1051 -1610
rect 1074 -1615 1075 -1610
rect 1079 -1615 1098 -1610
rect 130 -1626 134 -1623
rect 192 -1626 196 -1623
rect 130 -1630 162 -1626
rect 170 -1630 196 -1626
rect 933 -1622 937 -1616
rect 983 -1621 987 -1615
rect 1033 -1621 1037 -1615
rect 1080 -1621 1084 -1615
rect 90 -1648 94 -1645
rect 82 -1662 86 -1658
rect 130 -1662 134 -1630
rect 76 -1663 104 -1662
rect 76 -1667 96 -1663
rect 101 -1666 104 -1663
rect 109 -1666 134 -1662
rect 76 -1668 101 -1667
rect 941 -1686 945 -1672
rect 991 -1685 995 -1671
rect 1041 -1685 1045 -1671
rect 1088 -1685 1092 -1671
rect -278 -1719 -255 -1715
rect -274 -1721 -255 -1719
rect -278 -1730 -274 -1725
rect -259 -1730 -255 -1721
rect -242 -1726 -218 -1725
rect -242 -1730 -226 -1726
rect -222 -1730 -218 -1726
rect -242 -1732 -218 -1730
rect -236 -1737 -232 -1732
rect -267 -1758 -263 -1750
rect -267 -1762 -255 -1758
rect -259 -1764 -255 -1762
rect -228 -1764 -224 -1757
rect 2238 -1752 2277 -1751
rect 2238 -1756 2250 -1752
rect 2254 -1756 2360 -1752
rect 2238 -1758 2258 -1756
rect 2240 -1763 2244 -1758
rect 2286 -1760 2291 -1756
rect -284 -1769 -266 -1765
rect -259 -1768 -235 -1764
rect -228 -1768 -218 -1764
rect -284 -1776 -277 -1772
rect -259 -1779 -255 -1768
rect -228 -1771 -224 -1768
rect -236 -1785 -232 -1781
rect 2286 -1766 2291 -1764
rect -242 -1786 -217 -1785
rect -242 -1790 -222 -1786
rect -242 -1791 -217 -1790
rect 2248 -1790 2252 -1783
rect 2287 -1768 2291 -1766
rect 2305 -1768 2309 -1756
rect 2232 -1794 2241 -1790
rect 2248 -1794 2269 -1790
rect 2248 -1797 2252 -1794
rect -278 -1803 -274 -1799
rect -278 -1807 -262 -1803
rect 2240 -1811 2244 -1807
rect 2234 -1812 2259 -1811
rect 2234 -1814 2254 -1812
rect 2234 -1817 2247 -1814
rect 2253 -1816 2254 -1814
rect 2253 -1817 2259 -1816
rect 2265 -1821 2269 -1794
rect 2331 -1762 2353 -1759
rect 2331 -1768 2335 -1762
rect 2349 -1768 2353 -1762
rect 2296 -1812 2300 -1808
rect 2331 -1812 2335 -1808
rect 2296 -1816 2335 -1812
rect 2356 -1765 2360 -1756
rect 2356 -1770 2357 -1765
rect 2340 -1814 2344 -1808
rect 2340 -1818 2357 -1814
rect 2265 -1825 2332 -1821
rect 2269 -1833 2342 -1829
rect 1402 -1840 1422 -1836
rect 1433 -1840 1464 -1836
rect 1476 -1840 1504 -1836
rect 1514 -1840 1535 -1836
rect 1551 -1838 1581 -1834
rect 1402 -1843 1406 -1840
rect 1440 -1843 1444 -1840
rect 1484 -1843 1488 -1840
rect 1522 -1843 1526 -1840
rect 1568 -1841 1572 -1838
rect 1396 -1847 1397 -1843
rect 1401 -1847 1406 -1843
rect 1434 -1847 1435 -1843
rect 1439 -1847 1444 -1843
rect 1478 -1847 1479 -1843
rect 1483 -1847 1488 -1843
rect 1516 -1847 1517 -1843
rect 1521 -1847 1526 -1843
rect 1562 -1845 1563 -1841
rect 1567 -1845 1572 -1841
rect 94 -1857 133 -1856
rect 94 -1861 106 -1857
rect 110 -1861 216 -1857
rect 94 -1863 114 -1861
rect 96 -1868 100 -1863
rect 142 -1865 147 -1861
rect 142 -1871 147 -1869
rect 104 -1895 108 -1888
rect 143 -1873 147 -1871
rect 161 -1873 165 -1861
rect 88 -1899 97 -1895
rect 104 -1899 125 -1895
rect 104 -1902 108 -1899
rect 96 -1916 100 -1912
rect 90 -1917 115 -1916
rect 90 -1919 110 -1917
rect 90 -1922 103 -1919
rect 109 -1921 110 -1919
rect 109 -1922 115 -1921
rect 121 -1926 125 -1899
rect 187 -1867 209 -1864
rect 187 -1873 191 -1867
rect 205 -1873 209 -1867
rect 152 -1917 156 -1913
rect 187 -1917 191 -1913
rect 152 -1921 191 -1917
rect 212 -1870 216 -1861
rect 869 -1858 873 -1850
rect 897 -1858 901 -1850
rect 924 -1858 928 -1850
rect 963 -1858 967 -1850
rect 991 -1858 995 -1850
rect 1018 -1858 1022 -1850
rect 1058 -1857 1062 -1849
rect 1086 -1857 1090 -1849
rect 1113 -1857 1117 -1849
rect 1149 -1857 1153 -1849
rect 1402 -1853 1406 -1847
rect 1440 -1853 1444 -1847
rect 1484 -1853 1488 -1847
rect 1522 -1853 1526 -1847
rect 1568 -1851 1572 -1845
rect 2238 -1844 2257 -1843
rect 2238 -1848 2249 -1844
rect 2253 -1848 2257 -1844
rect 2238 -1850 2257 -1848
rect 212 -1875 213 -1870
rect 196 -1919 200 -1913
rect 196 -1923 213 -1919
rect 121 -1930 188 -1926
rect 125 -1938 198 -1934
rect 94 -1949 113 -1948
rect 94 -1953 105 -1949
rect 109 -1953 113 -1949
rect 94 -1955 113 -1953
rect 95 -1960 99 -1955
rect 103 -1987 107 -1980
rect 125 -1987 129 -1938
rect 209 -1942 213 -1923
rect 175 -1946 213 -1942
rect 175 -1949 179 -1946
rect 86 -1991 96 -1987
rect 103 -1991 129 -1987
rect 165 -1953 187 -1949
rect 2239 -1855 2243 -1850
rect 2247 -1882 2251 -1875
rect 2269 -1882 2273 -1833
rect 2353 -1837 2357 -1818
rect 2319 -1841 2357 -1837
rect 2319 -1844 2323 -1841
rect 2230 -1886 2240 -1882
rect 2247 -1886 2273 -1882
rect 2309 -1848 2331 -1844
rect 2287 -1867 2291 -1864
rect 2349 -1867 2353 -1864
rect 2287 -1871 2319 -1867
rect 2327 -1871 2353 -1867
rect 2247 -1889 2251 -1886
rect 1410 -1911 1414 -1893
rect 1448 -1911 1452 -1893
rect 1492 -1911 1496 -1893
rect 1530 -1911 1534 -1893
rect 1576 -1909 1580 -1891
rect 2239 -1903 2243 -1899
rect 2287 -1903 2291 -1871
rect 2233 -1904 2261 -1903
rect 2233 -1908 2253 -1904
rect 2258 -1907 2261 -1904
rect 2266 -1907 2291 -1903
rect 2233 -1909 2258 -1908
rect 1402 -1940 1406 -1931
rect 1440 -1940 1444 -1931
rect 1484 -1940 1488 -1931
rect 1522 -1940 1526 -1931
rect 1568 -1938 1572 -1929
rect 1402 -1944 1422 -1940
rect 1433 -1944 1464 -1940
rect 1476 -1944 1504 -1940
rect 1514 -1944 1531 -1940
rect 1551 -1942 1577 -1938
rect 877 -1964 881 -1958
rect 905 -1964 909 -1958
rect 932 -1964 936 -1958
rect 971 -1964 975 -1958
rect 999 -1964 1003 -1958
rect 1026 -1964 1030 -1958
rect 1066 -1963 1070 -1957
rect 1094 -1963 1098 -1957
rect 1121 -1963 1125 -1957
rect 1157 -1963 1161 -1957
rect 143 -1972 147 -1969
rect 205 -1972 209 -1969
rect 143 -1976 175 -1972
rect 183 -1976 209 -1972
rect 103 -1994 107 -1991
rect 95 -2008 99 -2004
rect 143 -2008 147 -1976
rect 89 -2009 117 -2008
rect 89 -2013 109 -2009
rect 114 -2012 117 -2009
rect 122 -2012 147 -2008
rect 89 -2014 114 -2013
rect -276 -2069 -253 -2065
rect -272 -2071 -253 -2069
rect -276 -2080 -272 -2075
rect -257 -2080 -253 -2071
rect -240 -2076 -216 -2075
rect -240 -2080 -224 -2076
rect -220 -2080 -216 -2076
rect -240 -2082 -216 -2080
rect -234 -2087 -230 -2082
rect -265 -2108 -261 -2100
rect -265 -2112 -253 -2108
rect -257 -2114 -253 -2112
rect -226 -2114 -222 -2107
rect -282 -2119 -264 -2115
rect -257 -2118 -233 -2114
rect -226 -2118 -216 -2114
rect -282 -2126 -275 -2122
rect -257 -2129 -253 -2118
rect -226 -2121 -222 -2118
rect 2240 -2121 2279 -2120
rect 2240 -2125 2252 -2121
rect 2256 -2125 2362 -2121
rect 2240 -2127 2260 -2125
rect -234 -2135 -230 -2131
rect 2242 -2132 2246 -2127
rect 2288 -2129 2293 -2125
rect -240 -2136 -215 -2135
rect -240 -2140 -220 -2136
rect -240 -2141 -215 -2140
rect -276 -2153 -272 -2149
rect -276 -2157 -260 -2153
rect 86 -2149 125 -2148
rect 86 -2153 98 -2149
rect 102 -2153 208 -2149
rect 2288 -2135 2293 -2133
rect 86 -2155 106 -2153
rect 88 -2160 92 -2155
rect 134 -2157 139 -2153
rect 134 -2163 139 -2161
rect 96 -2187 100 -2180
rect 135 -2165 139 -2163
rect 153 -2165 157 -2153
rect 80 -2191 89 -2187
rect 96 -2191 117 -2187
rect 96 -2194 100 -2191
rect 88 -2208 92 -2204
rect 82 -2209 107 -2208
rect 82 -2211 102 -2209
rect 82 -2214 95 -2211
rect 101 -2213 102 -2211
rect 101 -2214 107 -2213
rect 113 -2218 117 -2191
rect 179 -2159 201 -2156
rect 179 -2165 183 -2159
rect 197 -2165 201 -2159
rect 144 -2209 148 -2205
rect 179 -2209 183 -2205
rect 144 -2213 183 -2209
rect 204 -2162 208 -2153
rect 204 -2167 205 -2162
rect 2250 -2159 2254 -2152
rect 2289 -2137 2293 -2135
rect 2307 -2137 2311 -2125
rect 2234 -2163 2243 -2159
rect 2250 -2163 2271 -2159
rect 2250 -2166 2254 -2163
rect 2242 -2180 2246 -2176
rect 2236 -2181 2261 -2180
rect 2236 -2183 2256 -2181
rect 2236 -2186 2249 -2183
rect 2255 -2185 2256 -2183
rect 2255 -2186 2261 -2185
rect 2267 -2190 2271 -2163
rect 2333 -2131 2355 -2128
rect 2333 -2137 2337 -2131
rect 2351 -2137 2355 -2131
rect 2298 -2181 2302 -2177
rect 2333 -2181 2337 -2177
rect 2298 -2185 2337 -2181
rect 2358 -2134 2362 -2125
rect 2358 -2139 2359 -2134
rect 2342 -2183 2346 -2177
rect 2342 -2187 2359 -2183
rect 2267 -2194 2334 -2190
rect 2271 -2202 2344 -2198
rect 188 -2211 192 -2205
rect 188 -2215 205 -2211
rect 113 -2222 180 -2218
rect 117 -2230 190 -2226
rect 86 -2241 105 -2240
rect 86 -2245 97 -2241
rect 101 -2245 105 -2241
rect 86 -2247 105 -2245
rect 87 -2252 91 -2247
rect 95 -2279 99 -2272
rect 117 -2279 121 -2230
rect 201 -2234 205 -2215
rect 2240 -2213 2259 -2212
rect 2240 -2217 2251 -2213
rect 2255 -2217 2259 -2213
rect 2240 -2219 2259 -2217
rect 167 -2238 205 -2234
rect 2241 -2224 2245 -2219
rect 167 -2241 171 -2238
rect 78 -2283 88 -2279
rect 95 -2283 121 -2279
rect 157 -2245 179 -2241
rect 2249 -2251 2253 -2244
rect 2271 -2251 2275 -2202
rect 2355 -2206 2359 -2187
rect 2321 -2210 2359 -2206
rect 2321 -2213 2325 -2210
rect 2232 -2255 2242 -2251
rect 2249 -2255 2275 -2251
rect 2311 -2217 2333 -2213
rect 2289 -2236 2293 -2233
rect 2351 -2236 2355 -2233
rect 2289 -2240 2321 -2236
rect 2329 -2240 2355 -2236
rect 2249 -2258 2253 -2255
rect 135 -2264 139 -2261
rect 197 -2264 201 -2261
rect 135 -2268 167 -2264
rect 175 -2268 201 -2264
rect 95 -2286 99 -2283
rect 87 -2300 91 -2296
rect 135 -2300 139 -2268
rect 2241 -2272 2245 -2268
rect 2289 -2272 2293 -2240
rect 2235 -2273 2263 -2272
rect 2235 -2277 2255 -2273
rect 2260 -2276 2263 -2273
rect 2268 -2276 2293 -2272
rect 2235 -2278 2260 -2277
rect 81 -2301 109 -2300
rect 81 -2305 101 -2301
rect 106 -2304 109 -2301
rect 114 -2304 139 -2300
rect 81 -2306 106 -2305
rect -268 -2361 -245 -2357
rect -264 -2363 -245 -2361
rect -268 -2372 -264 -2367
rect -249 -2372 -245 -2363
rect -232 -2368 -208 -2367
rect -232 -2372 -216 -2368
rect -212 -2372 -208 -2368
rect -232 -2374 -208 -2372
rect -226 -2379 -222 -2374
rect -257 -2400 -253 -2392
rect -257 -2404 -245 -2400
rect -249 -2406 -245 -2404
rect -218 -2406 -214 -2399
rect -274 -2411 -256 -2407
rect -249 -2410 -225 -2406
rect -218 -2410 -208 -2406
rect -274 -2418 -267 -2414
rect -249 -2421 -245 -2410
rect -218 -2413 -214 -2410
rect -226 -2427 -222 -2423
rect -232 -2428 -207 -2427
rect -232 -2432 -212 -2428
rect -232 -2433 -207 -2432
rect -268 -2445 -264 -2441
rect -268 -2449 -252 -2445
rect 87 -2452 126 -2451
rect 87 -2456 99 -2452
rect 103 -2456 209 -2452
rect 87 -2458 107 -2456
rect 89 -2463 93 -2458
rect 135 -2460 140 -2456
rect 135 -2466 140 -2464
rect 97 -2490 101 -2483
rect 136 -2468 140 -2466
rect 154 -2468 158 -2456
rect 81 -2494 90 -2490
rect 97 -2494 118 -2490
rect 97 -2497 101 -2494
rect 89 -2511 93 -2507
rect 83 -2512 108 -2511
rect 83 -2514 103 -2512
rect 83 -2517 96 -2514
rect 102 -2516 103 -2514
rect 102 -2517 108 -2516
rect 114 -2521 118 -2494
rect 180 -2462 202 -2459
rect 180 -2468 184 -2462
rect 198 -2468 202 -2462
rect 145 -2512 149 -2508
rect 180 -2512 184 -2508
rect 145 -2516 184 -2512
rect 205 -2465 209 -2456
rect 2255 -2454 2294 -2453
rect 2255 -2458 2267 -2454
rect 2271 -2458 2377 -2454
rect 2255 -2460 2275 -2458
rect 2257 -2465 2261 -2460
rect 2303 -2462 2308 -2458
rect 205 -2470 206 -2465
rect 2303 -2468 2308 -2466
rect 2265 -2492 2269 -2485
rect 2304 -2470 2308 -2468
rect 2322 -2470 2326 -2458
rect 2249 -2496 2258 -2492
rect 2265 -2496 2286 -2492
rect 2265 -2499 2269 -2496
rect 189 -2514 193 -2508
rect 2257 -2513 2261 -2509
rect 2251 -2514 2276 -2513
rect 189 -2518 206 -2514
rect 114 -2525 181 -2521
rect 118 -2533 191 -2529
rect 87 -2544 106 -2543
rect 87 -2548 98 -2544
rect 102 -2548 106 -2544
rect 87 -2550 106 -2548
rect 88 -2555 92 -2550
rect 96 -2582 100 -2575
rect 118 -2582 122 -2533
rect 202 -2537 206 -2518
rect 2251 -2516 2271 -2514
rect 2251 -2519 2264 -2516
rect 2270 -2518 2271 -2516
rect 2270 -2519 2276 -2518
rect 2282 -2523 2286 -2496
rect 2348 -2464 2370 -2461
rect 2348 -2470 2352 -2464
rect 2366 -2470 2370 -2464
rect 2313 -2514 2317 -2510
rect 2348 -2514 2352 -2510
rect 2313 -2518 2352 -2514
rect 2373 -2467 2377 -2458
rect 2373 -2472 2374 -2467
rect 2357 -2516 2361 -2510
rect 2357 -2520 2374 -2516
rect 2282 -2527 2349 -2523
rect 168 -2541 206 -2537
rect 2286 -2535 2359 -2531
rect 168 -2544 172 -2541
rect 79 -2586 89 -2582
rect 96 -2586 122 -2582
rect 158 -2548 180 -2544
rect 2255 -2546 2274 -2545
rect 2255 -2550 2266 -2546
rect 2270 -2550 2274 -2546
rect 2255 -2552 2274 -2550
rect 136 -2567 140 -2564
rect 198 -2567 202 -2564
rect 136 -2571 168 -2567
rect 176 -2571 202 -2567
rect 2256 -2557 2260 -2552
rect 96 -2589 100 -2586
rect 88 -2603 92 -2599
rect 136 -2603 140 -2571
rect 2264 -2584 2268 -2577
rect 2286 -2584 2290 -2535
rect 2370 -2539 2374 -2520
rect 2336 -2543 2374 -2539
rect 2336 -2546 2340 -2543
rect 2247 -2588 2257 -2584
rect 2264 -2588 2290 -2584
rect 2326 -2550 2348 -2546
rect 2304 -2569 2308 -2566
rect 2366 -2569 2370 -2566
rect 2304 -2573 2336 -2569
rect 2344 -2573 2370 -2569
rect 2264 -2591 2268 -2588
rect 82 -2604 110 -2603
rect 82 -2608 102 -2604
rect 107 -2607 110 -2604
rect 115 -2607 140 -2603
rect 2256 -2605 2260 -2601
rect 2304 -2605 2308 -2573
rect 2250 -2606 2278 -2605
rect 82 -2609 107 -2608
rect 2250 -2610 2270 -2606
rect 2275 -2609 2278 -2606
rect 2283 -2609 2308 -2605
rect 2250 -2611 2275 -2610
rect -280 -2727 -257 -2723
rect -276 -2729 -257 -2727
rect -280 -2738 -276 -2733
rect -261 -2738 -257 -2729
rect -244 -2734 -220 -2733
rect -244 -2738 -228 -2734
rect -224 -2738 -220 -2734
rect -244 -2740 -220 -2738
rect -238 -2745 -234 -2740
rect -269 -2766 -265 -2758
rect -269 -2770 -257 -2766
rect -261 -2772 -257 -2770
rect -230 -2772 -226 -2765
rect -286 -2777 -268 -2773
rect -261 -2776 -237 -2772
rect -230 -2776 -220 -2772
rect -286 -2784 -279 -2780
rect -261 -2787 -257 -2776
rect -230 -2779 -226 -2776
rect -238 -2793 -234 -2789
rect -244 -2794 -219 -2793
rect -244 -2798 -224 -2794
rect -244 -2799 -219 -2798
rect -280 -2811 -276 -2807
rect -280 -2815 -264 -2811
<< m2contact >>
rect 2229 -1477 2235 -1471
rect 69 -1554 75 -1548
rect 2227 -1569 2233 -1563
rect 67 -1646 73 -1640
rect 2226 -1795 2232 -1789
rect 82 -1900 88 -1894
rect 80 -1992 86 -1986
rect 2224 -1887 2230 -1881
rect 74 -2192 80 -2186
rect 2228 -2164 2234 -2158
rect 72 -2284 78 -2278
rect 2226 -2256 2232 -2250
rect 75 -2495 81 -2489
rect 2243 -2497 2249 -2491
rect 73 -2587 79 -2581
rect 2241 -2589 2247 -2583
<< pm12contact >>
rect 932 -1695 938 -1689
rect 982 -1694 988 -1688
rect 1032 -1694 1038 -1688
rect 1079 -1694 1085 -1688
rect 1402 -1908 1407 -1903
rect 1440 -1908 1445 -1903
rect 1484 -1908 1489 -1903
rect 1522 -1908 1527 -1903
rect 1568 -1906 1573 -1901
rect 869 -1970 874 -1965
rect 897 -1970 902 -1965
rect 924 -1970 929 -1965
rect 963 -1970 968 -1965
rect 991 -1970 996 -1965
rect 1018 -1970 1023 -1965
rect 1058 -1969 1063 -1964
rect 1086 -1969 1091 -1964
rect 1113 -1969 1118 -1964
rect 1149 -1969 1154 -1964
<< pnm12contact >>
rect 2289 -1499 2296 -1494
rect 129 -1576 136 -1571
rect 2301 -1522 2307 -1518
rect 141 -1599 147 -1595
rect 2286 -1817 2293 -1812
rect 142 -1922 149 -1917
rect 154 -1945 160 -1941
rect 2298 -1840 2304 -1836
rect 134 -2214 141 -2209
rect 2288 -2186 2295 -2181
rect 146 -2237 152 -2233
rect 2300 -2209 2306 -2205
rect 135 -2517 142 -2512
rect 147 -2540 153 -2536
rect 2303 -2519 2310 -2514
rect 2315 -2542 2321 -2538
<< metal2 >>
rect 2230 -1482 2234 -1477
rect 2230 -1486 2279 -1482
rect 2275 -1495 2279 -1486
rect 2275 -1499 2289 -1495
rect 2228 -1518 2284 -1516
rect 2228 -1520 2301 -1518
rect 70 -1559 74 -1554
rect 70 -1563 119 -1559
rect 2228 -1563 2232 -1520
rect 2280 -1522 2301 -1520
rect 2280 -1523 2284 -1522
rect 115 -1572 119 -1563
rect 2233 -1568 2234 -1564
rect 115 -1576 129 -1572
rect 68 -1595 124 -1593
rect 68 -1597 141 -1595
rect 68 -1640 72 -1597
rect 120 -1599 141 -1597
rect 120 -1600 124 -1599
rect 73 -1645 74 -1641
rect 922 -1695 932 -1689
rect 972 -1694 982 -1688
rect 1022 -1694 1032 -1688
rect 1069 -1694 1079 -1688
rect 2227 -1800 2231 -1795
rect 2227 -1804 2276 -1800
rect 2272 -1813 2276 -1804
rect 2272 -1817 2286 -1813
rect 2225 -1836 2281 -1834
rect 2225 -1838 2298 -1836
rect 2225 -1881 2229 -1838
rect 2277 -1840 2298 -1838
rect 2277 -1841 2281 -1840
rect 2230 -1886 2231 -1882
rect 83 -1905 87 -1900
rect 83 -1909 132 -1905
rect 1399 -1908 1402 -1903
rect 1437 -1908 1440 -1903
rect 1481 -1908 1484 -1903
rect 1519 -1908 1522 -1903
rect 1565 -1906 1568 -1901
rect 128 -1918 132 -1909
rect 128 -1922 142 -1918
rect 81 -1941 137 -1939
rect 81 -1943 154 -1941
rect 81 -1986 85 -1943
rect 133 -1945 154 -1943
rect 133 -1946 137 -1945
rect 865 -1970 869 -1965
rect 893 -1970 897 -1965
rect 920 -1970 924 -1965
rect 959 -1970 963 -1965
rect 987 -1970 991 -1965
rect 1014 -1970 1018 -1965
rect 1054 -1969 1058 -1964
rect 1082 -1969 1086 -1964
rect 1109 -1969 1113 -1964
rect 1145 -1969 1149 -1964
rect 86 -1991 87 -1987
rect 2229 -2169 2233 -2164
rect 2229 -2173 2278 -2169
rect 2274 -2182 2278 -2173
rect 2274 -2186 2288 -2182
rect 75 -2197 79 -2192
rect 75 -2201 124 -2197
rect 120 -2210 124 -2201
rect 2227 -2205 2283 -2203
rect 2227 -2207 2300 -2205
rect 120 -2214 134 -2210
rect 73 -2233 129 -2231
rect 73 -2235 146 -2233
rect 73 -2278 77 -2235
rect 125 -2237 146 -2235
rect 125 -2238 129 -2237
rect 2227 -2250 2231 -2207
rect 2279 -2209 2300 -2207
rect 2279 -2210 2283 -2209
rect 2232 -2255 2233 -2251
rect 78 -2283 79 -2279
rect 76 -2500 80 -2495
rect 76 -2504 125 -2500
rect 121 -2513 125 -2504
rect 2244 -2502 2248 -2497
rect 2244 -2506 2293 -2502
rect 121 -2517 135 -2513
rect 2289 -2515 2293 -2506
rect 2289 -2519 2303 -2515
rect 74 -2536 130 -2534
rect 74 -2538 147 -2536
rect 74 -2581 78 -2538
rect 126 -2540 147 -2538
rect 2242 -2538 2298 -2536
rect 2242 -2540 2315 -2538
rect 126 -2541 130 -2540
rect 79 -2586 80 -2582
rect 2242 -2583 2246 -2540
rect 2294 -2542 2315 -2540
rect 2294 -2543 2298 -2542
rect 2247 -2588 2248 -2584
<< m123contact >>
rect 2235 -1440 2241 -1433
rect 2250 -1501 2256 -1496
rect 75 -1517 81 -1510
rect 2236 -1532 2241 -1525
rect 90 -1578 96 -1573
rect 2264 -1590 2269 -1585
rect 76 -1609 81 -1602
rect 104 -1667 109 -1662
rect 2232 -1758 2238 -1751
rect 2247 -1819 2253 -1814
rect 88 -1863 94 -1856
rect 2233 -1850 2238 -1843
rect 2261 -1908 2266 -1903
rect 103 -1924 109 -1919
rect 89 -1955 94 -1948
rect 117 -2013 122 -2008
rect 2234 -2127 2240 -2120
rect 80 -2155 86 -2148
rect 2249 -2188 2255 -2183
rect 95 -2216 101 -2211
rect 81 -2247 86 -2240
rect 2235 -2219 2240 -2212
rect 2263 -2277 2268 -2272
rect 109 -2305 114 -2300
rect 81 -2458 87 -2451
rect 2249 -2460 2255 -2453
rect 96 -2519 102 -2514
rect 2264 -2521 2270 -2516
rect 82 -2550 87 -2543
rect 2250 -2552 2255 -2545
rect 110 -2608 115 -2603
rect 2278 -2610 2283 -2605
<< metal3 >>
rect 77 -1602 81 -1517
rect 2237 -1525 2241 -1440
rect 2252 -1496 2256 -1494
rect 2252 -1507 2256 -1501
rect 2252 -1511 2268 -1507
rect 92 -1573 96 -1571
rect 92 -1584 96 -1578
rect 92 -1588 108 -1584
rect 104 -1662 108 -1588
rect 2264 -1585 2268 -1511
rect 2234 -1843 2238 -1758
rect 2249 -1814 2253 -1812
rect 2249 -1825 2253 -1819
rect 2249 -1829 2265 -1825
rect 90 -1948 94 -1863
rect 2261 -1903 2265 -1829
rect 105 -1919 109 -1917
rect 105 -1930 109 -1924
rect 105 -1934 121 -1930
rect 117 -2008 121 -1934
rect 82 -2240 86 -2155
rect 97 -2211 101 -2209
rect 2236 -2212 2240 -2127
rect 2251 -2183 2255 -2181
rect 2251 -2194 2255 -2188
rect 2251 -2198 2267 -2194
rect 97 -2222 101 -2216
rect 97 -2226 113 -2222
rect 109 -2300 113 -2226
rect 2263 -2272 2267 -2198
rect 83 -2543 87 -2458
rect 98 -2514 102 -2512
rect 98 -2525 102 -2519
rect 98 -2529 114 -2525
rect 110 -2603 114 -2529
rect 2251 -2545 2255 -2460
rect 2266 -2516 2270 -2514
rect 2266 -2527 2270 -2521
rect 2266 -2531 2282 -2527
rect 2278 -2605 2282 -2531
<< labels >>
rlabel metal1 869 -1854 873 -1850 1 pdr1
rlabel metal2 865 -1970 869 -1965 2 prop_1
rlabel metal1 877 -1964 881 -1959 1 prop1_car0
rlabel metal1 897 -1855 901 -1850 1 prop1_car0
rlabel metal2 893 -1970 897 -1965 1 carry_0
rlabel metal1 905 -1964 909 -1959 1 clock_car0
rlabel metal1 924 -1855 928 -1850 1 clock_car0
rlabel metal2 920 -1970 924 -1965 1 clock_in
rlabel metal1 932 -1964 936 -1959 1 gnd!
rlabel metal1 963 -1855 967 -1850 1 pdr2
rlabel metal2 959 -1970 963 -1965 1 prop_2
rlabel metal1 971 -1964 975 -1959 1 pdr1
rlabel metal1 991 -1855 995 -1850 1 pdr1
rlabel metal2 987 -1970 991 -1965 1 gen_1
rlabel metal1 999 -1964 1003 -1959 1 clock_car0
rlabel metal1 1018 -1855 1022 -1850 1 pdr3
rlabel metal2 1014 -1970 1018 -1965 1 prop_3
rlabel metal1 1026 -1964 1030 -1959 1 pdr2
rlabel metal1 1058 -1854 1062 -1849 1 pdr2
rlabel metal2 1054 -1969 1058 -1964 1 gen_2
rlabel metal1 1066 -1963 1070 -1958 1 clock_car0
rlabel metal1 1086 -1854 1090 -1849 1 pdr4
rlabel metal2 1082 -1969 1086 -1964 1 prop_4
rlabel metal1 1094 -1963 1098 -1958 1 pdr3
rlabel metal1 1113 -1854 1117 -1849 1 pdr3
rlabel metal2 1109 -1969 1113 -1964 1 gen_3
rlabel metal1 1121 -1963 1125 -1958 1 clock_car0
rlabel metal1 1149 -1854 1153 -1849 1 pdr4
rlabel metal2 1145 -1969 1149 -1964 1 gen_4
rlabel metal1 1157 -1963 1161 -1958 7 clock_car0
rlabel metal1 933 -1607 937 -1602 5 vdd!
rlabel metal1 983 -1606 987 -1601 5 vdd!
rlabel metal1 1033 -1606 1037 -1601 5 vdd!
rlabel metal1 1080 -1606 1084 -1601 5 vdd!
rlabel metal2 922 -1695 928 -1689 2 clock_in
rlabel metal2 972 -1694 978 -1688 1 clock_in
rlabel metal2 1022 -1694 1028 -1688 1 clock_in
rlabel metal2 1069 -1694 1074 -1688 1 clock_in
rlabel metal1 941 -1686 945 -1681 1 pdr1
rlabel metal1 991 -1685 995 -1681 1 pdr2
rlabel metal1 1041 -1685 1045 -1681 1 pdr3
rlabel metal1 1088 -1685 1092 -1681 1 pdr4
rlabel metal1 1527 -1944 1531 -1940 1 gnd!
rlabel metal1 1523 -1840 1528 -1836 5 vdd!
rlabel metal2 1399 -1908 1402 -1903 1 pdr1
rlabel metal2 1437 -1908 1440 -1903 1 pdr2
rlabel metal2 1481 -1908 1484 -1903 1 pdr3
rlabel metal2 1519 -1908 1522 -1903 1 pdr4
rlabel metal1 1410 -1908 1414 -1903 1 c1
rlabel metal1 1448 -1908 1452 -1903 1 c2
rlabel metal1 1492 -1908 1496 -1903 1 c3
rlabel metal1 1530 -1908 1534 -1903 1 c4
rlabel metal1 1573 -1942 1577 -1938 1 gnd!
rlabel metal1 1569 -1838 1574 -1834 5 vdd!
rlabel metal2 1565 -1906 1568 -1901 1 clk_org
rlabel metal1 1576 -1906 1580 -1901 1 clock_in
rlabel metal1 1402 -1840 1406 -1836 5 vdd!
rlabel metal1 1440 -1840 1444 -1836 5 vdd!
rlabel metal1 1484 -1840 1488 -1836 5 vdd!
rlabel metal1 1488 -1944 1492 -1940 1 gnd!
rlabel metal1 1451 -1944 1455 -1940 1 gnd!
rlabel metal1 1411 -1944 1415 -1940 1 gnd!
rlabel metal1 150 -1513 150 -1513 5 vdd
rlabel metal1 162 -1628 162 -1628 1 gnd
rlabel m123contact 80 -1607 80 -1607 5 vdd
rlabel metal1 83 -1664 83 -1664 1 gnd
rlabel metal1 81 -1515 81 -1515 5 vdd
rlabel metal1 84 -1572 84 -1572 1 gnd
rlabel metal1 163 -1859 163 -1859 5 vdd
rlabel metal1 175 -1974 175 -1974 1 gnd
rlabel m123contact 93 -1953 93 -1953 5 vdd
rlabel metal1 96 -2010 96 -2010 1 gnd
rlabel metal1 94 -1861 94 -1861 5 vdd
rlabel metal1 97 -1918 97 -1918 1 gnd
rlabel metal1 155 -2151 155 -2151 5 vdd
rlabel metal1 167 -2266 167 -2266 1 gnd
rlabel m123contact 85 -2245 85 -2245 5 vdd
rlabel metal1 88 -2302 88 -2302 1 gnd
rlabel metal1 86 -2153 86 -2153 5 vdd
rlabel metal1 89 -2210 89 -2210 1 gnd
rlabel metal1 156 -2454 156 -2454 5 vdd
rlabel metal1 168 -2569 168 -2569 1 gnd
rlabel m123contact 86 -2548 86 -2548 5 vdd
rlabel metal1 89 -2605 89 -2605 1 gnd
rlabel metal1 87 -2456 87 -2456 5 vdd
rlabel metal1 90 -2513 90 -2513 1 gnd
rlabel metal1 2310 -1436 2310 -1436 5 vdd
rlabel metal1 2322 -1551 2322 -1551 1 gnd
rlabel m123contact 2240 -1530 2240 -1530 5 vdd
rlabel metal1 2243 -1587 2243 -1587 1 gnd
rlabel metal1 2241 -1438 2241 -1438 5 vdd
rlabel metal1 2244 -1495 2244 -1495 1 gnd
rlabel metal1 2307 -1754 2307 -1754 5 vdd
rlabel metal1 2319 -1869 2319 -1869 1 gnd
rlabel m123contact 2237 -1848 2237 -1848 5 vdd
rlabel metal1 2240 -1905 2240 -1905 1 gnd
rlabel metal1 2238 -1756 2238 -1756 5 vdd
rlabel metal1 2241 -1813 2241 -1813 1 gnd
rlabel metal1 2309 -2123 2309 -2123 5 vdd
rlabel metal1 2321 -2238 2321 -2238 1 gnd
rlabel m123contact 2239 -2217 2239 -2217 5 vdd
rlabel metal1 2242 -2274 2242 -2274 1 gnd
rlabel metal1 2240 -2125 2240 -2125 5 vdd
rlabel metal1 2243 -2182 2243 -2182 1 gnd
rlabel metal1 2324 -2456 2324 -2456 5 vdd
rlabel metal1 2336 -2571 2336 -2571 1 gnd
rlabel m123contact 2254 -2550 2254 -2550 5 vdd
rlabel metal1 2257 -2607 2257 -2607 1 gnd
rlabel metal1 2255 -2458 2255 -2458 5 vdd
rlabel metal1 2258 -2515 2258 -2515 1 gnd
rlabel metal1 -268 -1718 -268 -1718 5 vdd
rlabel metal1 -267 -1805 -267 -1805 1 gnd
rlabel metal1 -235 -1787 -235 -1787 1 gnd
rlabel metal1 -238 -1730 -238 -1730 5 vdd
rlabel metal1 -266 -2068 -266 -2068 5 vdd
rlabel metal1 -265 -2155 -265 -2155 1 gnd
rlabel metal1 -233 -2137 -233 -2137 1 gnd
rlabel metal1 -236 -2080 -236 -2080 5 vdd
rlabel metal1 -258 -2360 -258 -2360 5 vdd
rlabel metal1 -257 -2447 -257 -2447 1 gnd
rlabel metal1 -225 -2429 -225 -2429 1 gnd
rlabel metal1 -228 -2372 -228 -2372 5 vdd
rlabel metal1 -270 -2726 -270 -2726 5 vdd
rlabel metal1 -269 -2813 -269 -2813 1 gnd
rlabel metal1 -237 -2795 -237 -2795 1 gnd
rlabel metal1 -240 -2738 -240 -2738 5 vdd
rlabel metal2 70 -1616 70 -1616 1 q_b1
rlabel metal2 71 -1560 71 -1560 1 q_a1
rlabel metal1 198 -1585 198 -1585 1 prop_1
rlabel metal1 -283 -1767 -283 -1767 3 q_a1
rlabel metal1 -281 -1774 -281 -1774 3 q_b1
rlabel metal2 84 -1905 84 -1905 1 q_a2
rlabel metal2 84 -1965 84 -1965 1 q_b2
rlabel metal1 211 -1935 211 -1935 1 prop_2
rlabel metal1 -219 -1767 -219 -1767 1 gen_1
rlabel metal1 -280 -2118 -280 -2118 1 q_a2
rlabel metal1 -280 -2125 -280 -2125 1 q_b2
rlabel metal1 -217 -2116 -217 -2116 1 gen_2
rlabel metal2 76 -2196 76 -2196 1 q_a3
rlabel metal2 75 -2235 75 -2235 1 q_b3
rlabel metal1 204 -2227 204 -2227 1 prop_3
rlabel metal1 -273 -2410 -273 -2410 1 q_b3
rlabel metal1 -271 -2417 -271 -2417 1 q_a3
rlabel metal1 -210 -2408 -210 -2408 1 gen_3
rlabel metal2 78 -2500 78 -2500 1 q_b4
rlabel metal1 204 -2524 204 -2524 1 prop_4
rlabel metal2 75 -2555 75 -2555 1 q_a4
rlabel metal1 -285 -2775 -285 -2775 3 q_a4
rlabel metal1 -285 -2781 -285 -2781 3 q_b4
rlabel metal1 -222 -2774 -222 -2774 1 gen_4
rlabel m2contact 2231 -1473 2231 -1473 1 carry_0
rlabel m2contact 2228 -1567 2228 -1567 1 prop_1
rlabel metal1 2358 -1505 2358 -1505 1 s1
rlabel metal1 2355 -1830 2355 -1830 1 s2
rlabel metal1 2358 -2196 2358 -2196 1 s3
rlabel metal1 2372 -2528 2372 -2528 1 s4
rlabel m2contact 2230 -1792 2230 -1792 1 c1
rlabel m2contact 2230 -2162 2230 -2162 1 c2
rlabel m2contact 2247 -2495 2247 -2495 1 c3
rlabel m2contact 2244 -2587 2244 -2587 1 prop_4
rlabel m2contact 2229 -2253 2229 -2253 1 prop_3
rlabel m2contact 2227 -1884 2227 -1884 1 prop_2
<< end >>
