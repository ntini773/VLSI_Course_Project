magic
tech scmos
timestamp 1732005981
<< nwell >>
rect 485 140 509 180
rect 529 170 566 172
rect 529 115 567 170
rect 573 115 616 167
rect 484 48 508 88
<< ntransistor >>
rect 496 122 498 132
rect 543 65 545 85
rect 553 65 555 85
rect 587 65 589 85
rect 597 65 599 85
rect 495 30 497 40
<< ptransistor >>
rect 496 146 498 166
rect 543 121 545 161
rect 553 121 555 161
rect 587 121 589 161
rect 597 121 599 161
rect 495 54 497 74
<< ndiffusion >>
rect 495 122 496 132
rect 498 122 499 132
rect 542 65 543 85
rect 545 65 553 85
rect 555 65 556 85
rect 586 65 587 85
rect 589 65 597 85
rect 599 65 600 85
rect 494 30 495 40
rect 497 30 498 40
<< pdiffusion >>
rect 495 146 496 166
rect 498 146 499 166
rect 542 121 543 161
rect 545 121 547 161
rect 551 121 553 161
rect 555 121 556 161
rect 586 121 587 161
rect 589 121 591 161
rect 595 121 597 161
rect 599 121 600 161
rect 494 54 495 74
rect 497 54 498 74
<< ndcontact >>
rect 491 122 495 132
rect 499 122 503 132
rect 538 65 542 85
rect 556 65 560 85
rect 582 65 586 85
rect 600 65 604 85
rect 490 30 494 40
rect 498 30 502 40
<< pdcontact >>
rect 491 146 495 166
rect 499 146 503 166
rect 538 121 542 161
rect 547 121 551 161
rect 556 121 560 161
rect 582 121 586 161
rect 591 121 595 161
rect 600 121 604 161
rect 490 54 494 74
rect 498 54 502 74
<< psubstratepcontact >>
rect 505 113 510 117
rect 570 58 578 62
rect 504 21 509 25
<< nsubstratencontact >>
rect 501 173 505 177
rect 537 165 543 169
rect 608 159 613 164
rect 500 81 504 85
<< polysilicon >>
rect 496 166 498 170
rect 543 161 545 164
rect 553 161 555 164
rect 587 161 589 164
rect 597 161 599 164
rect 496 132 498 146
rect 496 119 498 122
rect 543 117 545 121
rect 544 112 545 117
rect 543 85 545 112
rect 553 93 555 121
rect 553 85 555 89
rect 587 85 589 121
rect 597 85 599 121
rect 495 74 497 78
rect 543 62 545 65
rect 553 62 555 65
rect 587 62 589 65
rect 597 62 599 65
rect 495 40 497 54
rect 495 27 497 30
<< polycontact >>
rect 492 135 496 139
rect 583 104 587 108
rect 593 96 597 100
rect 491 43 495 47
<< metal1 >>
rect 489 177 528 178
rect 489 173 501 177
rect 505 173 611 177
rect 489 171 509 173
rect 491 166 495 171
rect 537 169 542 173
rect 537 163 542 165
rect 499 139 503 146
rect 538 161 542 163
rect 556 161 560 173
rect 483 135 492 139
rect 499 135 520 139
rect 499 132 503 135
rect 491 118 495 122
rect 485 117 510 118
rect 485 115 505 117
rect 485 112 498 115
rect 504 113 505 115
rect 504 112 510 113
rect 516 108 520 135
rect 582 167 604 170
rect 582 161 586 167
rect 600 161 604 167
rect 547 117 551 121
rect 582 117 586 121
rect 547 113 586 117
rect 607 164 611 173
rect 607 159 608 164
rect 591 115 595 121
rect 591 111 608 115
rect 516 104 583 108
rect 520 96 593 100
rect 489 85 508 86
rect 489 81 500 85
rect 504 81 508 85
rect 489 79 508 81
rect 490 74 494 79
rect 498 47 502 54
rect 520 47 524 96
rect 604 92 608 111
rect 570 88 608 92
rect 570 85 574 88
rect 481 43 491 47
rect 498 43 524 47
rect 560 81 582 85
rect 538 62 542 65
rect 600 62 604 65
rect 538 58 570 62
rect 578 58 604 62
rect 498 40 502 43
rect 490 26 494 30
rect 538 26 542 58
rect 484 25 512 26
rect 484 21 504 25
rect 509 22 512 25
rect 517 22 542 26
rect 484 20 509 21
<< m2contact >>
rect 477 134 483 140
rect 475 42 481 48
<< pnm12contact >>
rect 537 112 544 117
rect 549 89 555 93
<< metal2 >>
rect 478 129 482 134
rect 478 125 527 129
rect 523 116 527 125
rect 523 112 537 116
rect 476 93 532 95
rect 476 91 549 93
rect 476 48 480 91
rect 528 89 549 91
rect 528 88 532 89
rect 481 43 482 47
<< m123contact >>
rect 483 171 489 178
rect 498 110 504 115
rect 484 79 489 86
rect 512 21 517 26
<< metal3 >>
rect 485 86 489 171
rect 500 115 504 117
rect 500 104 504 110
rect 500 100 516 104
rect 512 26 516 100
<< labels >>
rlabel metal1 558 175 558 175 5 vdd
rlabel metal1 606 106 606 106 7 out
rlabel metal1 570 60 570 60 1 gnd
rlabel m123contact 488 81 488 81 5 vdd
rlabel metal1 491 24 491 24 1 gnd
rlabel metal1 506 45 506 45 1 out
rlabel metal1 489 173 489 173 5 vdd
rlabel metal1 492 116 492 116 1 gnd
rlabel metal1 507 137 507 137 1 out
<< end >>
