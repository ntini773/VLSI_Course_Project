magic
tech scmos
timestamp 1731944955
<< nwell >>
rect 852 143 876 205
rect 882 143 906 205
rect 912 143 936 205
rect 945 143 969 205
<< ntransistor >>
rect 854 16 856 116
rect 882 16 884 116
rect 909 16 911 116
rect 948 16 950 116
rect 976 16 978 116
rect 1003 16 1005 116
rect 1043 17 1045 117
rect 1071 17 1073 117
rect 1098 17 1100 117
rect 1134 17 1136 117
<< ptransistor >>
rect 863 149 865 199
rect 893 149 895 199
rect 923 149 925 199
rect 956 149 958 199
<< ndiffusion >>
rect 853 16 854 116
rect 856 16 857 116
rect 881 16 882 116
rect 884 16 885 116
rect 908 16 909 116
rect 911 16 912 116
rect 947 16 948 116
rect 950 16 951 116
rect 975 16 976 116
rect 978 16 979 116
rect 1002 16 1003 116
rect 1005 16 1006 116
rect 1042 17 1043 117
rect 1045 17 1046 117
rect 1070 17 1071 117
rect 1073 17 1074 117
rect 1097 17 1098 117
rect 1100 17 1101 117
rect 1133 17 1134 117
rect 1136 17 1137 117
<< pdiffusion >>
rect 862 149 863 199
rect 865 149 866 199
rect 892 149 893 199
rect 895 149 896 199
rect 922 149 923 199
rect 925 149 926 199
rect 955 149 956 199
rect 958 149 959 199
<< ndcontact >>
rect 849 16 853 116
rect 857 16 861 116
rect 877 16 881 116
rect 885 16 889 116
rect 904 16 908 116
rect 912 16 916 116
rect 943 16 947 116
rect 951 16 955 116
rect 971 16 975 116
rect 979 16 983 116
rect 998 16 1002 116
rect 1006 16 1010 116
rect 1038 17 1042 117
rect 1046 17 1050 117
rect 1066 17 1070 117
rect 1074 17 1078 117
rect 1093 17 1097 117
rect 1101 17 1105 117
rect 1129 17 1133 117
rect 1137 17 1141 117
<< pdcontact >>
rect 858 149 862 199
rect 866 149 870 199
rect 888 149 892 199
rect 896 149 900 199
rect 918 149 922 199
rect 926 149 930 199
rect 951 149 955 199
rect 959 149 963 199
<< nsubstratencontact >>
rect 853 205 857 209
rect 883 205 887 209
rect 913 205 917 209
rect 946 205 950 209
<< polysilicon >>
rect 863 199 865 202
rect 893 199 895 202
rect 923 199 925 202
rect 956 199 958 202
rect 863 134 865 149
rect 893 134 895 149
rect 923 134 925 149
rect 956 134 958 149
rect 854 116 856 119
rect 882 116 884 119
rect 909 116 911 119
rect 948 116 950 119
rect 976 116 978 119
rect 1003 116 1005 119
rect 1043 117 1045 120
rect 1071 117 1073 120
rect 1098 117 1100 120
rect 1134 117 1136 120
rect 854 4 856 16
rect 882 4 884 16
rect 909 4 911 16
rect 948 4 950 16
rect 976 4 978 16
rect 1003 4 1005 16
rect 1043 5 1045 17
rect 1071 5 1073 17
rect 1098 5 1100 17
rect 1134 5 1136 17
<< metal1 >>
rect 858 209 862 212
rect 888 209 892 212
rect 918 209 922 212
rect 951 209 955 212
rect 852 205 853 209
rect 857 205 862 209
rect 882 205 883 209
rect 887 205 892 209
rect 912 205 913 209
rect 917 205 922 209
rect 945 205 946 209
rect 950 205 955 209
rect 858 199 862 205
rect 888 199 892 205
rect 918 199 922 205
rect 951 199 955 205
rect 867 139 870 149
rect 897 139 900 149
rect 927 139 930 149
rect 960 139 963 149
rect 849 116 853 124
rect 877 116 881 124
rect 904 116 908 124
rect 943 116 947 124
rect 971 116 975 124
rect 998 116 1002 124
rect 1038 117 1042 125
rect 1066 117 1070 125
rect 1093 117 1097 125
rect 1129 117 1133 125
rect 857 10 861 16
rect 885 10 889 16
rect 912 10 916 16
rect 951 10 955 16
rect 979 10 983 16
rect 1006 10 1010 16
rect 1046 11 1050 17
rect 1074 11 1078 17
rect 1101 11 1105 17
rect 1137 11 1141 17
<< pm12contact >>
rect 858 134 863 139
rect 888 134 893 139
rect 918 134 923 139
rect 951 134 956 139
rect 849 4 854 9
rect 877 4 882 9
rect 904 4 909 9
rect 943 4 948 9
rect 971 4 976 9
rect 998 4 1003 9
rect 1038 5 1043 10
rect 1066 5 1071 10
rect 1093 5 1098 10
rect 1129 5 1134 10
<< metal2 >>
rect 855 134 858 139
rect 885 134 888 139
rect 915 134 918 139
rect 948 134 951 139
rect 845 4 849 9
rect 873 4 877 9
rect 900 4 904 9
rect 939 4 943 9
rect 967 4 971 9
rect 994 4 998 9
rect 1034 5 1038 10
rect 1062 5 1066 10
rect 1089 5 1093 10
rect 1125 5 1129 10
<< labels >>
rlabel metal1 858 209 862 212 5 vdd!
rlabel metal1 888 209 892 212 5 vdd!
rlabel metal1 918 209 922 212 5 vdd!
rlabel metal2 855 134 858 139 2 clock_in
rlabel metal2 885 134 888 139 1 clock_in
rlabel metal2 915 134 918 139 1 clock_in
rlabel metal2 948 134 951 139 1 clock_in
rlabel metal1 867 139 870 142 1 pdr1
rlabel metal1 897 139 900 142 1 pdr2
rlabel metal1 927 139 930 142 1 pdr3
rlabel metal1 960 139 963 142 1 pdr4
rlabel metal1 849 120 853 124 1 pdr1
rlabel metal2 845 4 849 9 2 prop_1
rlabel metal1 857 10 861 15 1 prop1_car0
rlabel metal1 877 119 881 124 1 prop1_car0
rlabel metal2 873 4 877 9 1 carry_0
rlabel metal1 885 10 889 15 1 clock_car0
rlabel metal1 904 119 908 124 1 clock_car0
rlabel metal2 900 4 904 9 1 clock_in
rlabel metal1 912 10 916 15 1 gnd!
rlabel metal1 943 119 947 124 1 pdr2
rlabel metal2 939 4 943 9 1 prop_2
rlabel metal1 951 10 955 15 1 pdr1
rlabel metal1 971 119 975 124 1 pdr1
rlabel metal2 967 4 971 9 1 gen_1
rlabel metal1 979 10 983 15 1 clock_car0
rlabel metal1 998 119 1002 124 1 pdr3
rlabel metal2 994 4 998 9 1 prop_3
rlabel metal1 1006 10 1010 15 1 pdr2
rlabel metal1 1038 120 1042 125 1 pdr2
rlabel metal2 1034 5 1038 10 1 gen_2
rlabel metal1 1046 11 1050 16 1 clock_car0
rlabel metal1 1066 120 1070 125 1 pdr4
rlabel metal2 1062 5 1066 10 1 prop_4
rlabel metal1 1074 11 1078 16 1 pdr3
rlabel metal1 1093 120 1097 125 1 pdr3
rlabel metal2 1089 5 1093 10 1 gen_3
rlabel metal1 1101 11 1105 16 1 clock_car0
rlabel metal1 1129 120 1133 125 1 pdr4
rlabel metal2 1125 5 1129 10 1 gen_4
rlabel metal1 1137 11 1141 16 7 clock_car0
<< end >>
