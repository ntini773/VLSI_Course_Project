magic
tech scmos
timestamp 1732006825
<< nwell >>
rect 218 120 242 160
rect 262 150 299 152
rect 262 95 300 150
rect 306 95 349 147
rect 217 28 241 68
<< ntransistor >>
rect 229 102 231 112
rect 276 45 278 65
rect 286 45 288 65
rect 320 45 322 65
rect 330 45 332 65
rect 228 10 230 20
<< ptransistor >>
rect 229 126 231 146
rect 276 101 278 141
rect 286 101 288 141
rect 320 101 322 141
rect 330 101 332 141
rect 228 34 230 54
<< ndiffusion >>
rect 228 102 229 112
rect 231 102 232 112
rect 275 45 276 65
rect 278 45 286 65
rect 288 45 289 65
rect 319 45 320 65
rect 322 45 330 65
rect 332 45 333 65
rect 227 10 228 20
rect 230 10 231 20
<< pdiffusion >>
rect 228 126 229 146
rect 231 126 232 146
rect 275 101 276 141
rect 278 101 280 141
rect 284 101 286 141
rect 288 101 289 141
rect 319 101 320 141
rect 322 101 324 141
rect 328 101 330 141
rect 332 101 333 141
rect 227 34 228 54
rect 230 34 231 54
<< ndcontact >>
rect 224 102 228 112
rect 232 102 236 112
rect 271 45 275 65
rect 289 45 293 65
rect 315 45 319 65
rect 333 45 337 65
rect 223 10 227 20
rect 231 10 235 20
<< pdcontact >>
rect 224 126 228 146
rect 232 126 236 146
rect 271 101 275 141
rect 280 101 284 141
rect 289 101 293 141
rect 315 101 319 141
rect 324 101 328 141
rect 333 101 337 141
rect 223 34 227 54
rect 231 34 235 54
<< psubstratepcontact >>
rect 238 93 243 97
rect 303 38 311 42
rect 237 1 242 5
<< nsubstratencontact >>
rect 234 153 238 157
rect 270 145 276 149
rect 341 139 346 144
rect 233 61 237 65
<< polysilicon >>
rect 229 146 231 150
rect 276 141 278 144
rect 286 141 288 144
rect 320 141 322 144
rect 330 141 332 144
rect 229 112 231 126
rect 229 99 231 102
rect 276 97 278 101
rect 277 92 278 97
rect 276 65 278 92
rect 286 73 288 101
rect 286 65 288 69
rect 320 65 322 101
rect 330 65 332 101
rect 228 54 230 58
rect 276 42 278 45
rect 286 42 288 45
rect 320 42 322 45
rect 330 42 332 45
rect 228 20 230 34
rect 228 7 230 10
<< polycontact >>
rect 225 115 229 119
rect 316 84 320 88
rect 326 76 330 80
rect 224 23 228 27
<< metal1 >>
rect 222 157 261 158
rect 222 153 234 157
rect 238 153 344 157
rect 222 151 242 153
rect 224 146 228 151
rect 270 149 275 153
rect 270 143 275 145
rect 232 119 236 126
rect 271 141 275 143
rect 289 141 293 153
rect 216 115 225 119
rect 232 115 253 119
rect 232 112 236 115
rect 224 98 228 102
rect 218 97 243 98
rect 218 95 238 97
rect 218 92 231 95
rect 237 93 238 95
rect 237 92 243 93
rect 249 88 253 115
rect 315 147 337 150
rect 315 141 319 147
rect 333 141 337 147
rect 280 97 284 101
rect 315 97 319 101
rect 280 93 319 97
rect 340 144 344 153
rect 340 139 341 144
rect 324 95 328 101
rect 324 91 341 95
rect 249 84 316 88
rect 253 76 326 80
rect 222 65 241 66
rect 222 61 233 65
rect 237 61 241 65
rect 222 59 241 61
rect 223 54 227 59
rect 231 27 235 34
rect 253 27 257 76
rect 337 72 341 91
rect 303 68 341 72
rect 303 65 307 68
rect 214 23 224 27
rect 231 23 257 27
rect 293 61 315 65
rect 271 42 275 45
rect 333 42 337 45
rect 271 38 303 42
rect 311 38 337 42
rect 231 20 235 23
rect 223 6 227 10
rect 271 6 275 38
rect 217 5 245 6
rect 217 1 237 5
rect 242 2 245 5
rect 250 2 275 6
rect 217 0 242 1
<< m2contact >>
rect 210 114 216 120
rect 208 22 214 28
<< pnm12contact >>
rect 270 92 277 97
rect 282 69 288 73
<< metal2 >>
rect 211 109 215 114
rect 211 105 260 109
rect 256 96 260 105
rect 256 92 270 96
rect 209 73 265 75
rect 209 71 282 73
rect 209 28 213 71
rect 261 69 282 71
rect 261 68 265 69
rect 214 23 215 27
<< m123contact >>
rect 216 151 222 158
rect 231 90 237 95
rect 217 59 222 66
rect 245 1 250 6
<< metal3 >>
rect 218 66 222 151
rect 233 95 237 97
rect 233 84 237 90
rect 233 80 249 84
rect 245 6 249 80
<< labels >>
rlabel metal1 291 155 291 155 5 vdd
rlabel metal1 303 40 303 40 1 gnd
rlabel m123contact 221 61 221 61 5 vdd
rlabel metal1 224 4 224 4 1 gnd
rlabel metal1 222 153 222 153 5 vdd
rlabel metal1 225 96 225 96 1 gnd
<< end >>
