magic
tech scmos
timestamp 1732005398
<< nwell >>
rect -11 -14 25 26
rect 31 -21 55 19
<< ntransistor >>
rect 0 -57 2 -37
rect 11 -57 13 -37
rect 42 -39 44 -29
<< ptransistor >>
rect 0 -8 2 12
rect 11 -8 13 12
rect 42 -15 44 5
<< ndiffusion >>
rect -1 -57 0 -37
rect 2 -57 11 -37
rect 13 -57 14 -37
rect 41 -39 42 -29
rect 44 -39 45 -29
<< pdiffusion >>
rect -1 -8 0 12
rect 2 -8 6 12
rect 10 -8 11 12
rect 13 -8 14 12
rect 41 -15 42 5
rect 44 -15 45 5
<< ndcontact >>
rect -5 -57 -1 -37
rect 14 -57 18 -37
rect 37 -39 41 -29
rect 45 -39 49 -29
<< pdcontact >>
rect -5 -8 -1 12
rect 6 -8 10 12
rect 14 -8 18 12
rect 37 -15 41 5
rect 45 -15 49 5
<< psubstratepcontact >>
rect 51 -48 56 -44
<< nsubstratencontact >>
rect -5 17 -1 23
rect 47 12 51 16
<< polysilicon >>
rect 0 12 2 15
rect 11 12 13 15
rect 42 5 44 9
rect 0 -37 2 -8
rect 11 -37 13 -8
rect 42 -29 44 -15
rect 42 -42 44 -39
rect 0 -60 2 -57
rect 11 -60 13 -57
<< polycontact >>
rect -4 -34 0 -30
rect 7 -27 11 -23
rect 38 -26 42 -22
<< metal1 >>
rect -5 23 18 27
rect -1 21 18 23
rect -5 12 -1 17
rect 14 12 18 21
rect 31 16 55 17
rect 31 12 47 16
rect 51 12 55 16
rect 31 10 55 12
rect 37 5 41 10
rect 6 -16 10 -8
rect 6 -20 18 -16
rect 14 -22 18 -20
rect 45 -22 49 -15
rect -11 -27 7 -23
rect 14 -26 38 -22
rect 45 -26 55 -22
rect -11 -34 -4 -30
rect 14 -37 18 -26
rect 45 -29 49 -26
rect 37 -43 41 -39
rect 31 -44 56 -43
rect 31 -48 51 -44
rect 31 -49 56 -48
rect -5 -61 -1 -57
rect -5 -65 11 -61
<< labels >>
rlabel metal1 5 24 5 24 5 vdd
rlabel metal1 6 -63 6 -63 1 gnd
rlabel metal1 38 -45 38 -45 1 gnd
rlabel metal1 35 12 35 12 5 vdd
<< end >>
