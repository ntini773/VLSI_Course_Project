magic
tech scmos
timestamp 1731655617
<< nwell >>
rect -9 -25 17 14
rect 47 -25 73 14
rect 107 -25 133 14
rect -9 -96 17 -57
<< ntransistor >>
rect 58 -72 60 -62
rect 122 -74 124 -64
rect 2 -143 4 -133
rect 50 -134 52 -124
rect 108 -131 110 -121
<< ptransistor >>
rect 3 -13 5 7
rect 59 -13 61 7
rect 119 -13 121 7
rect 4 -88 6 -68
<< ndiffusion >>
rect 57 -72 58 -62
rect 60 -72 61 -62
rect 121 -74 122 -64
rect 124 -74 125 -64
rect 1 -143 2 -133
rect 4 -143 5 -133
rect 49 -134 50 -124
rect 52 -134 53 -124
rect 107 -131 108 -121
rect 110 -131 111 -121
<< pdiffusion >>
rect 2 -13 3 7
rect 5 -13 6 7
rect 58 -13 59 7
rect 61 -13 62 7
rect 118 -13 119 7
rect 121 -13 122 7
rect 3 -88 4 -68
rect 6 -88 7 -68
<< ndcontact >>
rect 53 -72 57 -62
rect 61 -72 65 -62
rect 117 -74 121 -64
rect 125 -74 129 -64
rect -3 -143 1 -133
rect 5 -143 9 -133
rect 45 -134 49 -124
rect 53 -134 57 -124
rect 103 -131 107 -121
rect 111 -131 115 -121
<< pdcontact >>
rect -2 -13 2 7
rect 6 -13 10 7
rect 54 -13 58 7
rect 62 -13 66 7
rect 114 -13 118 7
rect 122 -13 126 7
rect -1 -88 3 -68
rect 7 -88 11 -68
<< polysilicon >>
rect 3 7 5 19
rect 59 7 61 16
rect 119 7 121 17
rect 3 -31 5 -13
rect 59 -32 61 -13
rect 119 -40 121 -13
rect 58 -62 60 -59
rect 4 -68 6 -62
rect 122 -64 124 -59
rect 58 -78 60 -72
rect 4 -102 6 -88
rect 122 -89 124 -74
rect 108 -121 110 -117
rect 50 -124 52 -121
rect 2 -133 4 -130
rect 50 -143 52 -134
rect 2 -146 4 -143
rect 108 -145 110 -131
<< polycontact >>
rect 1 -36 5 -31
rect 57 -36 61 -32
rect 117 -44 121 -40
rect 56 -82 60 -78
rect 119 -95 124 -89
rect 2 -107 6 -102
rect 0 -130 4 -126
rect 48 -147 52 -143
rect 105 -150 110 -145
<< metal1 >>
rect -10 21 136 27
rect -2 7 2 21
rect 54 7 58 21
rect 114 7 118 21
rect 6 -25 10 -13
rect 6 -28 24 -25
rect -15 -36 1 -31
rect -15 -91 -12 -36
rect 20 -51 24 -28
rect 62 -26 66 -13
rect 62 -29 77 -26
rect 38 -36 57 -32
rect 73 -40 77 -29
rect 122 -28 126 -13
rect 193 -28 196 -25
rect 122 -32 196 -28
rect 242 -29 265 -25
rect 73 -44 117 -40
rect 73 -45 77 -44
rect -1 -54 24 -51
rect 53 -50 77 -45
rect -1 -68 3 -54
rect 53 -62 57 -50
rect 61 -75 71 -72
rect -24 -95 -12 -91
rect 7 -92 11 -88
rect 47 -82 56 -78
rect 47 -92 50 -82
rect 7 -95 50 -92
rect -24 -126 -21 -95
rect 7 -96 11 -95
rect -15 -107 2 -102
rect 20 -108 23 -95
rect 12 -112 23 -108
rect 67 -109 71 -75
rect -24 -130 0 -126
rect -3 -153 1 -143
rect 12 -143 16 -112
rect 45 -113 71 -109
rect 45 -124 49 -113
rect 53 -135 57 -134
rect 53 -138 64 -135
rect 5 -148 16 -143
rect 36 -147 48 -143
rect 61 -153 64 -138
rect 87 -145 91 -44
rect 149 -49 154 -32
rect 117 -54 154 -49
rect 117 -64 121 -54
rect 149 -65 154 -54
rect 125 -77 129 -74
rect 125 -80 152 -77
rect 100 -95 119 -89
rect 148 -107 152 -80
rect 103 -111 152 -107
rect 103 -121 107 -111
rect 111 -137 115 -131
rect 111 -140 135 -137
rect 87 -150 105 -145
rect 129 -153 135 -140
rect -13 -157 135 -153
use inv  inv_0
timestamp 1731617906
transform 1 0 203 0 1 -7
box -7 -55 39 29
<< labels >>
rlabel metal1 -11 -33 -11 -33 3 d
rlabel metal1 4 24 4 24 5 vdd
rlabel metal1 22 -29 22 -29 7 c
rlabel metal1 -9 -105 -9 -105 1 clk
rlabel metal1 16 -111 16 -111 1 x
rlabel metal1 0 -155 0 -155 1 gnd
rlabel metal1 73 -28 73 -27 1 y
rlabel metal1 39 -145 39 -145 1 clk_2
rlabel metal1 103 -90 103 -90 1 clk_3
rlabel metal1 150 -98 150 -98 1 b
rlabel metal1 70 -97 70 -97 1 a
rlabel metal1 46 -34 46 -34 1 clk_1
<< end >>
