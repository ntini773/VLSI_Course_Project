magic
tech scmos
timestamp 1731964643
<< nwell >>
rect 309 601 342 648
rect 361 607 427 649
rect 112 508 145 555
rect 178 512 210 550
rect 306 307 339 354
rect 358 313 424 355
rect 885 313 909 375
rect 935 314 959 376
rect 985 314 1009 376
rect 1032 314 1056 376
rect 1777 374 1810 421
rect 1829 380 1895 422
rect 85 249 118 296
rect 151 253 183 291
rect 1792 164 1825 211
rect 1844 170 1910 212
rect 301 86 334 133
rect 353 92 419 134
rect 1354 92 1378 144
rect 1392 92 1416 144
rect 1436 92 1460 144
rect 1474 92 1498 144
rect 1520 94 1544 146
rect 66 -60 99 -13
rect 132 -56 164 -18
rect 1797 -65 1830 -18
rect 1849 -59 1915 -17
rect 314 -247 347 -200
rect 366 -241 432 -199
rect 1797 -256 1830 -209
rect 1849 -250 1915 -208
rect 71 -434 104 -387
rect 137 -430 169 -392
<< ntransistor >>
rect 325 583 327 593
rect 374 580 376 590
rect 408 580 410 590
rect 128 490 130 500
rect 192 481 194 491
rect 183 429 185 439
rect 322 289 324 299
rect 1793 356 1795 366
rect 1842 353 1844 363
rect 1876 353 1878 363
rect 371 286 373 296
rect 405 286 407 296
rect 101 231 103 241
rect 165 222 167 232
rect 156 170 158 180
rect 1808 146 1810 156
rect 1857 143 1859 153
rect 1891 143 1893 153
rect 317 68 319 78
rect 366 65 368 75
rect 400 65 402 75
rect 832 33 834 133
rect 860 33 862 133
rect 887 33 889 133
rect 926 33 928 133
rect 954 33 956 133
rect 981 33 983 133
rect 1021 34 1023 134
rect 1049 34 1051 134
rect 1076 34 1078 134
rect 1112 34 1114 134
rect 1365 60 1367 80
rect 1403 60 1405 80
rect 1447 60 1449 80
rect 1485 60 1487 80
rect 1531 62 1533 82
rect 82 -78 84 -68
rect 146 -87 148 -77
rect 1813 -83 1815 -73
rect 1862 -86 1864 -76
rect 1896 -86 1898 -76
rect 137 -139 139 -129
rect 330 -265 332 -255
rect 379 -268 381 -258
rect 413 -268 415 -258
rect 1813 -274 1815 -264
rect 1862 -277 1864 -267
rect 1896 -277 1898 -267
rect 87 -452 89 -442
rect 151 -461 153 -451
rect 142 -513 144 -503
<< ptransistor >>
rect 325 613 327 633
rect 374 621 376 641
rect 408 621 410 641
rect 128 520 130 540
rect 192 523 194 543
rect 1793 386 1795 406
rect 1842 394 1844 414
rect 1876 394 1878 414
rect 322 319 324 339
rect 371 327 373 347
rect 405 327 407 347
rect 896 319 898 369
rect 946 320 948 370
rect 996 320 998 370
rect 1043 320 1045 370
rect 101 261 103 281
rect 165 264 167 284
rect 1808 176 1810 196
rect 1857 184 1859 204
rect 1891 184 1893 204
rect 317 98 319 118
rect 366 106 368 126
rect 400 106 402 126
rect 1365 98 1367 138
rect 1403 98 1405 138
rect 1447 98 1449 138
rect 1485 98 1487 138
rect 1531 100 1533 140
rect 82 -48 84 -28
rect 146 -45 148 -25
rect 1813 -53 1815 -33
rect 1862 -45 1864 -25
rect 1896 -45 1898 -25
rect 330 -235 332 -215
rect 379 -227 381 -207
rect 413 -227 415 -207
rect 1813 -244 1815 -224
rect 1862 -236 1864 -216
rect 1896 -236 1898 -216
rect 87 -422 89 -402
rect 151 -419 153 -399
<< ndiffusion >>
rect 324 583 325 593
rect 327 583 328 593
rect 373 580 374 590
rect 376 580 377 590
rect 407 580 408 590
rect 410 580 411 590
rect 127 490 128 500
rect 130 490 131 500
rect 191 481 192 491
rect 194 481 195 491
rect 182 429 183 439
rect 185 429 186 439
rect 321 289 322 299
rect 324 289 325 299
rect 1792 356 1793 366
rect 1795 356 1796 366
rect 1841 353 1842 363
rect 1844 353 1845 363
rect 1875 353 1876 363
rect 1878 353 1879 363
rect 370 286 371 296
rect 373 286 374 296
rect 404 286 405 296
rect 407 286 408 296
rect 100 231 101 241
rect 103 231 104 241
rect 164 222 165 232
rect 167 222 168 232
rect 155 170 156 180
rect 158 170 159 180
rect 1807 146 1808 156
rect 1810 146 1811 156
rect 1856 143 1857 153
rect 1859 143 1860 153
rect 1890 143 1891 153
rect 1893 143 1894 153
rect 316 68 317 78
rect 319 68 320 78
rect 365 65 366 75
rect 368 65 369 75
rect 399 65 400 75
rect 402 65 403 75
rect 831 33 832 133
rect 834 33 835 133
rect 859 33 860 133
rect 862 33 863 133
rect 886 33 887 133
rect 889 33 890 133
rect 925 33 926 133
rect 928 33 929 133
rect 953 33 954 133
rect 956 33 957 133
rect 980 33 981 133
rect 983 33 984 133
rect 1020 34 1021 134
rect 1023 34 1024 134
rect 1048 34 1049 134
rect 1051 34 1052 134
rect 1075 34 1076 134
rect 1078 34 1079 134
rect 1111 34 1112 134
rect 1114 34 1115 134
rect 1364 60 1365 80
rect 1367 60 1368 80
rect 1402 60 1403 80
rect 1405 60 1406 80
rect 1446 60 1447 80
rect 1449 60 1450 80
rect 1484 60 1485 80
rect 1487 60 1488 80
rect 1530 62 1531 82
rect 1533 62 1534 82
rect 81 -78 82 -68
rect 84 -78 85 -68
rect 145 -87 146 -77
rect 148 -87 149 -77
rect 1812 -83 1813 -73
rect 1815 -83 1816 -73
rect 1861 -86 1862 -76
rect 1864 -86 1865 -76
rect 1895 -86 1896 -76
rect 1898 -86 1899 -76
rect 136 -139 137 -129
rect 139 -139 140 -129
rect 329 -265 330 -255
rect 332 -265 333 -255
rect 378 -268 379 -258
rect 381 -268 382 -258
rect 412 -268 413 -258
rect 415 -268 416 -258
rect 1812 -274 1813 -264
rect 1815 -274 1816 -264
rect 1861 -277 1862 -267
rect 1864 -277 1865 -267
rect 1895 -277 1896 -267
rect 1898 -277 1899 -267
rect 86 -452 87 -442
rect 89 -452 90 -442
rect 150 -461 151 -451
rect 153 -461 154 -451
rect 141 -513 142 -503
rect 144 -513 145 -503
<< pdiffusion >>
rect 324 613 325 633
rect 327 613 328 633
rect 373 621 374 641
rect 376 621 377 641
rect 407 621 408 641
rect 410 621 411 641
rect 127 520 128 540
rect 130 520 131 540
rect 191 523 192 543
rect 194 523 195 543
rect 1792 386 1793 406
rect 1795 386 1796 406
rect 1841 394 1842 414
rect 1844 394 1845 414
rect 1875 394 1876 414
rect 1878 394 1879 414
rect 321 319 322 339
rect 324 319 325 339
rect 370 327 371 347
rect 373 327 374 347
rect 404 327 405 347
rect 407 327 408 347
rect 895 319 896 369
rect 898 319 899 369
rect 945 320 946 370
rect 948 320 949 370
rect 995 320 996 370
rect 998 320 999 370
rect 1042 320 1043 370
rect 1045 320 1046 370
rect 100 261 101 281
rect 103 261 104 281
rect 164 264 165 284
rect 167 264 168 284
rect 1807 176 1808 196
rect 1810 176 1811 196
rect 1856 184 1857 204
rect 1859 184 1860 204
rect 1890 184 1891 204
rect 1893 184 1894 204
rect 316 98 317 118
rect 319 98 320 118
rect 365 106 366 126
rect 368 106 369 126
rect 399 106 400 126
rect 402 106 403 126
rect 1364 98 1365 138
rect 1367 98 1368 138
rect 1402 98 1403 138
rect 1405 98 1406 138
rect 1446 98 1447 138
rect 1449 98 1450 138
rect 1484 98 1485 138
rect 1487 98 1488 138
rect 1530 100 1531 140
rect 1533 100 1534 140
rect 81 -48 82 -28
rect 84 -48 85 -28
rect 145 -45 146 -25
rect 148 -45 149 -25
rect 1812 -53 1813 -33
rect 1815 -53 1816 -33
rect 1861 -45 1862 -25
rect 1864 -45 1865 -25
rect 1895 -45 1896 -25
rect 1898 -45 1899 -25
rect 329 -235 330 -215
rect 332 -235 333 -215
rect 378 -227 379 -207
rect 381 -227 382 -207
rect 412 -227 413 -207
rect 415 -227 416 -207
rect 1812 -244 1813 -224
rect 1815 -244 1816 -224
rect 1861 -236 1862 -216
rect 1864 -236 1865 -216
rect 1895 -236 1896 -216
rect 1898 -236 1899 -216
rect 86 -422 87 -402
rect 89 -422 90 -402
rect 150 -419 151 -399
rect 153 -419 154 -399
<< ndcontact >>
rect 320 583 324 593
rect 328 583 332 593
rect 369 580 373 590
rect 377 580 381 590
rect 403 580 407 590
rect 411 580 415 590
rect 123 490 127 500
rect 131 490 135 500
rect 187 481 191 491
rect 195 481 199 491
rect 178 429 182 439
rect 186 429 190 439
rect 317 289 321 299
rect 325 289 329 299
rect 1788 356 1792 366
rect 1796 356 1800 366
rect 1837 353 1841 363
rect 1845 353 1849 363
rect 1871 353 1875 363
rect 1879 353 1883 363
rect 366 286 370 296
rect 374 286 378 296
rect 400 286 404 296
rect 408 286 412 296
rect 96 231 100 241
rect 104 231 108 241
rect 160 222 164 232
rect 168 222 172 232
rect 151 170 155 180
rect 159 170 163 180
rect 1803 146 1807 156
rect 1811 146 1815 156
rect 1852 143 1856 153
rect 1860 143 1864 153
rect 1886 143 1890 153
rect 1894 143 1898 153
rect 312 68 316 78
rect 320 68 324 78
rect 361 65 365 75
rect 369 65 373 75
rect 395 65 399 75
rect 403 65 407 75
rect 827 33 831 133
rect 835 33 839 133
rect 855 33 859 133
rect 863 33 867 133
rect 882 33 886 133
rect 890 33 894 133
rect 921 33 925 133
rect 929 33 933 133
rect 949 33 953 133
rect 957 33 961 133
rect 976 33 980 133
rect 984 33 988 133
rect 1016 34 1020 134
rect 1024 34 1028 134
rect 1044 34 1048 134
rect 1052 34 1056 134
rect 1071 34 1075 134
rect 1079 34 1083 134
rect 1107 34 1111 134
rect 1115 34 1119 134
rect 1360 60 1364 80
rect 1368 60 1372 80
rect 1398 60 1402 80
rect 1406 60 1410 80
rect 1442 60 1446 80
rect 1450 60 1454 80
rect 1480 60 1484 80
rect 1488 60 1492 80
rect 1526 62 1530 82
rect 1534 62 1538 82
rect 77 -78 81 -68
rect 85 -78 89 -68
rect 141 -87 145 -77
rect 149 -87 153 -77
rect 1808 -83 1812 -73
rect 1816 -83 1820 -73
rect 1857 -86 1861 -76
rect 1865 -86 1869 -76
rect 1891 -86 1895 -76
rect 1899 -86 1903 -76
rect 132 -139 136 -129
rect 140 -139 144 -129
rect 325 -265 329 -255
rect 333 -265 337 -255
rect 374 -268 378 -258
rect 382 -268 386 -258
rect 408 -268 412 -258
rect 416 -268 420 -258
rect 1808 -274 1812 -264
rect 1816 -274 1820 -264
rect 1857 -277 1861 -267
rect 1865 -277 1869 -267
rect 1891 -277 1895 -267
rect 1899 -277 1903 -267
rect 82 -452 86 -442
rect 90 -452 94 -442
rect 146 -461 150 -451
rect 154 -461 158 -451
rect 137 -513 141 -503
rect 145 -513 149 -503
<< pdcontact >>
rect 320 613 324 633
rect 328 613 332 633
rect 369 621 373 641
rect 377 621 381 641
rect 403 621 407 641
rect 411 621 415 641
rect 123 520 127 540
rect 131 520 135 540
rect 187 523 191 543
rect 195 523 199 543
rect 1788 386 1792 406
rect 1796 386 1800 406
rect 1837 394 1841 414
rect 1845 394 1849 414
rect 1871 394 1875 414
rect 1879 394 1883 414
rect 317 319 321 339
rect 325 319 329 339
rect 366 327 370 347
rect 374 327 378 347
rect 400 327 404 347
rect 408 327 412 347
rect 891 319 895 369
rect 899 319 903 369
rect 941 320 945 370
rect 949 320 953 370
rect 991 320 995 370
rect 999 320 1003 370
rect 1038 320 1042 370
rect 1046 320 1050 370
rect 96 261 100 281
rect 104 261 108 281
rect 160 264 164 284
rect 168 264 172 284
rect 1803 176 1807 196
rect 1811 176 1815 196
rect 1852 184 1856 204
rect 1860 184 1864 204
rect 1886 184 1890 204
rect 1894 184 1898 204
rect 312 98 316 118
rect 320 98 324 118
rect 361 106 365 126
rect 369 106 373 126
rect 395 106 399 126
rect 403 106 407 126
rect 1360 98 1364 138
rect 1368 98 1372 138
rect 1398 98 1402 138
rect 1406 98 1410 138
rect 1442 98 1446 138
rect 1450 98 1454 138
rect 1480 98 1484 138
rect 1488 98 1492 138
rect 1526 100 1530 140
rect 1534 100 1538 140
rect 77 -48 81 -28
rect 85 -48 89 -28
rect 141 -45 145 -25
rect 149 -45 153 -25
rect 1808 -53 1812 -33
rect 1816 -53 1820 -33
rect 1857 -45 1861 -25
rect 1865 -45 1869 -25
rect 1891 -45 1895 -25
rect 1899 -45 1903 -25
rect 325 -235 329 -215
rect 333 -235 337 -215
rect 374 -227 378 -207
rect 382 -227 386 -207
rect 408 -227 412 -207
rect 416 -227 420 -207
rect 1808 -244 1812 -224
rect 1816 -244 1820 -224
rect 1857 -236 1861 -216
rect 1865 -236 1869 -216
rect 1891 -236 1895 -216
rect 1899 -236 1903 -216
rect 82 -422 86 -402
rect 90 -422 94 -402
rect 146 -419 150 -399
rect 154 -419 158 -399
<< nsubstratencontact >>
rect 886 375 890 380
rect 936 376 940 381
rect 986 376 990 381
rect 1033 376 1037 381
rect 1355 144 1359 148
rect 1393 144 1397 148
rect 1437 144 1441 148
rect 1475 144 1479 148
rect 1521 146 1525 150
<< polysilicon >>
rect 325 633 327 642
rect 374 641 376 648
rect 408 641 410 645
rect 325 593 327 613
rect 374 606 376 621
rect 374 590 376 593
rect 408 590 410 621
rect 325 580 327 583
rect 374 561 376 580
rect 408 577 410 580
rect 128 540 130 549
rect 192 543 194 553
rect 128 500 130 520
rect 192 508 194 523
rect 192 491 194 496
rect 128 487 130 490
rect 192 476 194 481
rect 183 439 185 460
rect 183 422 185 429
rect 1793 406 1795 415
rect 1842 414 1844 421
rect 1876 414 1878 418
rect 896 369 898 372
rect 946 370 948 373
rect 996 370 998 373
rect 1043 370 1045 373
rect 322 339 324 348
rect 371 347 373 354
rect 405 347 407 351
rect 322 299 324 319
rect 371 312 373 327
rect 101 281 103 290
rect 165 284 167 294
rect 371 296 373 299
rect 405 296 407 327
rect 1793 366 1795 386
rect 1842 379 1844 394
rect 1842 363 1844 366
rect 1876 363 1878 394
rect 1793 353 1795 356
rect 1842 334 1844 353
rect 1876 350 1878 353
rect 896 296 898 319
rect 946 297 948 320
rect 996 297 998 320
rect 1043 297 1045 320
rect 322 286 324 289
rect 371 267 373 286
rect 405 283 407 286
rect 101 241 103 261
rect 165 249 167 264
rect 165 232 167 237
rect 101 228 103 231
rect 165 217 167 222
rect 156 180 158 201
rect 1808 196 1810 205
rect 1857 204 1859 211
rect 1891 204 1893 208
rect 156 163 158 170
rect 1808 156 1810 176
rect 1857 169 1859 184
rect 1857 153 1859 156
rect 1891 153 1893 184
rect 1808 143 1810 146
rect 1365 138 1367 141
rect 1403 138 1405 141
rect 1447 138 1449 141
rect 1485 138 1487 141
rect 1531 140 1533 143
rect 832 133 834 136
rect 860 133 862 136
rect 887 133 889 136
rect 926 133 928 136
rect 954 133 956 136
rect 981 133 983 136
rect 1021 134 1023 137
rect 1049 134 1051 137
rect 1076 134 1078 137
rect 1112 134 1114 137
rect 317 118 319 127
rect 366 126 368 133
rect 400 126 402 130
rect 317 78 319 98
rect 366 91 368 106
rect 366 75 368 78
rect 400 75 402 106
rect 317 65 319 68
rect 366 46 368 65
rect 400 62 402 65
rect 1857 124 1859 143
rect 1891 140 1893 143
rect 1365 80 1367 98
rect 1403 80 1405 98
rect 1447 80 1449 98
rect 1485 80 1487 98
rect 1531 82 1533 100
rect 1365 56 1367 60
rect 1403 56 1405 60
rect 1447 56 1449 60
rect 1485 56 1487 60
rect 1531 58 1533 62
rect 832 21 834 33
rect 860 21 862 33
rect 887 21 889 33
rect 926 21 928 33
rect 954 21 956 33
rect 981 21 983 33
rect 1021 22 1023 34
rect 1049 22 1051 34
rect 1076 22 1078 34
rect 1112 22 1114 34
rect 82 -28 84 -19
rect 146 -25 148 -15
rect 1813 -33 1815 -24
rect 1862 -25 1864 -18
rect 1896 -25 1898 -21
rect 82 -68 84 -48
rect 146 -60 148 -45
rect 146 -77 148 -72
rect 1813 -73 1815 -53
rect 1862 -60 1864 -45
rect 82 -81 84 -78
rect 1862 -76 1864 -73
rect 1896 -76 1898 -45
rect 1813 -86 1815 -83
rect 146 -92 148 -87
rect 1862 -105 1864 -86
rect 1896 -89 1898 -86
rect 137 -129 139 -108
rect 137 -146 139 -139
rect 330 -215 332 -206
rect 379 -207 381 -200
rect 413 -207 415 -203
rect 1813 -224 1815 -215
rect 1862 -216 1864 -209
rect 1896 -216 1898 -212
rect 330 -255 332 -235
rect 379 -242 381 -227
rect 379 -258 381 -255
rect 413 -258 415 -227
rect 330 -268 332 -265
rect 1813 -264 1815 -244
rect 1862 -251 1864 -236
rect 379 -287 381 -268
rect 413 -271 415 -268
rect 1862 -267 1864 -264
rect 1896 -267 1898 -236
rect 1813 -277 1815 -274
rect 1862 -296 1864 -277
rect 1896 -280 1898 -277
rect 87 -402 89 -393
rect 151 -399 153 -389
rect 87 -442 89 -422
rect 151 -434 153 -419
rect 151 -451 153 -446
rect 87 -455 89 -452
rect 151 -466 153 -461
rect 142 -503 144 -482
rect 142 -520 144 -513
<< polycontact >>
rect 376 644 380 648
rect 321 596 325 600
rect 404 597 408 601
rect 376 561 381 566
rect 188 553 194 560
rect 124 503 128 507
rect 188 469 194 476
rect 181 460 185 464
rect 1844 417 1848 421
rect 373 350 377 354
rect 318 302 322 306
rect 161 294 167 301
rect 401 303 405 307
rect 1789 369 1793 373
rect 1872 370 1876 374
rect 1844 334 1849 339
rect 373 267 378 272
rect 97 244 101 248
rect 161 210 167 217
rect 154 201 158 205
rect 1859 207 1863 211
rect 1804 159 1808 163
rect 1887 160 1891 164
rect 368 129 372 133
rect 313 81 317 85
rect 396 82 400 86
rect 368 46 373 51
rect 1859 124 1864 129
rect 142 -15 148 -8
rect 1864 -22 1868 -18
rect 78 -65 82 -61
rect 1809 -70 1813 -66
rect 1892 -69 1896 -65
rect 142 -99 148 -92
rect 135 -108 139 -104
rect 1864 -105 1869 -100
rect 381 -204 385 -200
rect 1864 -213 1868 -209
rect 326 -252 330 -248
rect 409 -251 413 -247
rect 1809 -261 1813 -257
rect 1892 -260 1896 -256
rect 381 -287 386 -282
rect 1864 -296 1869 -291
rect 147 -389 153 -382
rect 83 -439 87 -435
rect 147 -473 153 -466
rect 140 -482 144 -478
<< metal1 >>
rect 352 671 359 680
rect 386 662 393 678
rect 294 658 393 662
rect 294 600 303 658
rect 309 648 352 655
rect 386 648 393 658
rect 320 633 324 648
rect 380 644 407 648
rect 403 641 407 644
rect 294 596 321 600
rect 328 599 332 613
rect 369 602 373 621
rect 328 595 355 599
rect 328 593 332 595
rect 320 578 324 583
rect 309 571 345 578
rect 89 565 163 570
rect 89 438 95 565
rect 112 555 145 562
rect 159 560 163 565
rect 123 540 127 555
rect 159 553 188 560
rect 350 557 355 595
rect 369 590 373 596
rect 369 574 373 580
rect 377 590 381 621
rect 411 602 415 621
rect 397 597 404 601
rect 411 596 435 602
rect 411 590 415 596
rect 398 584 403 590
rect 377 573 381 580
rect 411 573 415 580
rect 377 569 415 573
rect 381 561 385 566
rect 101 507 108 510
rect 101 503 124 507
rect 131 506 135 520
rect 159 507 166 553
rect 350 549 391 557
rect 158 506 166 507
rect 101 456 106 503
rect 131 502 166 506
rect 187 504 191 523
rect 131 500 135 502
rect 170 498 191 504
rect 187 491 191 498
rect 123 485 127 490
rect 112 478 148 485
rect 368 525 373 537
rect 195 505 199 523
rect 195 499 230 505
rect 195 491 199 499
rect 162 469 188 476
rect 162 456 169 469
rect 101 450 169 456
rect 173 460 181 464
rect 173 446 176 460
rect 224 456 230 499
rect 170 442 176 446
rect 186 450 230 456
rect 170 438 173 442
rect 186 439 190 450
rect 89 434 173 438
rect 1820 444 1827 453
rect 1854 435 1861 451
rect 1762 431 1861 435
rect 178 416 182 429
rect 166 411 202 416
rect 349 377 356 386
rect 383 368 390 384
rect 891 380 895 389
rect 941 381 945 390
rect 991 381 995 390
rect 1038 381 1042 390
rect 885 375 886 380
rect 890 375 909 380
rect 935 376 936 381
rect 940 376 959 381
rect 985 376 986 381
rect 990 376 1009 381
rect 1032 376 1033 381
rect 1037 376 1056 381
rect 291 364 390 368
rect 62 306 136 311
rect 62 179 68 306
rect 85 296 118 303
rect 132 301 136 306
rect 291 306 300 364
rect 306 354 349 361
rect 383 354 390 364
rect 891 369 895 375
rect 941 370 945 376
rect 991 370 995 376
rect 1038 370 1042 376
rect 1762 373 1771 431
rect 1777 421 1820 428
rect 1854 421 1861 431
rect 1788 406 1792 421
rect 1848 417 1875 421
rect 1871 414 1875 417
rect 317 339 321 354
rect 377 350 404 354
rect 400 347 404 350
rect 291 302 318 306
rect 325 305 329 319
rect 366 308 370 327
rect 325 301 352 305
rect 96 281 100 296
rect 132 294 161 301
rect 325 299 329 301
rect 74 248 81 251
rect 74 244 97 248
rect 104 247 108 261
rect 132 248 139 294
rect 317 284 321 289
rect 131 247 139 248
rect 74 197 79 244
rect 104 243 139 247
rect 160 245 164 264
rect 104 241 108 243
rect 143 239 164 245
rect 160 232 164 239
rect 96 226 100 231
rect 85 219 121 226
rect 306 277 342 284
rect 168 246 172 264
rect 347 263 352 301
rect 366 296 370 302
rect 366 280 370 286
rect 374 296 378 327
rect 408 308 412 327
rect 1762 369 1789 373
rect 1796 372 1800 386
rect 1837 375 1841 394
rect 1796 368 1823 372
rect 1796 366 1800 368
rect 1788 351 1792 356
rect 1777 344 1813 351
rect 1818 330 1823 368
rect 1837 363 1841 369
rect 1837 347 1841 353
rect 1845 363 1849 394
rect 1879 375 1883 394
rect 1865 370 1872 374
rect 1879 369 1903 375
rect 1879 363 1883 369
rect 1866 357 1871 363
rect 1845 346 1849 353
rect 1879 346 1883 353
rect 1845 342 1883 346
rect 1849 334 1853 339
rect 1818 322 1859 330
rect 394 303 401 307
rect 408 302 432 308
rect 899 305 903 319
rect 949 306 953 320
rect 999 306 1003 320
rect 1046 306 1050 320
rect 408 296 412 302
rect 1836 298 1841 310
rect 395 290 400 296
rect 374 279 378 286
rect 408 279 412 286
rect 374 275 412 279
rect 378 267 382 272
rect 347 255 388 263
rect 168 240 203 246
rect 168 232 172 240
rect 135 210 161 217
rect 135 197 142 210
rect 74 191 142 197
rect 146 201 154 205
rect 146 187 149 201
rect 197 197 203 240
rect 365 231 370 243
rect 1835 234 1842 243
rect 1869 225 1876 241
rect 143 183 149 187
rect 159 191 203 197
rect 1777 221 1876 225
rect 143 179 146 183
rect 159 180 163 191
rect 62 175 146 179
rect 151 157 155 170
rect 139 152 175 157
rect 344 156 351 165
rect 1777 163 1786 221
rect 1792 211 1835 218
rect 1869 211 1876 221
rect 1803 196 1807 211
rect 1863 207 1890 211
rect 1886 204 1890 207
rect 378 147 385 163
rect 1777 159 1804 163
rect 1811 162 1815 176
rect 1852 165 1856 184
rect 1811 158 1838 162
rect 1360 151 1380 155
rect 1391 151 1422 155
rect 1434 151 1462 155
rect 1472 151 1493 155
rect 1509 153 1539 157
rect 1811 156 1815 158
rect 1360 148 1364 151
rect 1398 148 1402 151
rect 1442 148 1446 151
rect 1480 148 1484 151
rect 1526 150 1530 153
rect 286 143 385 147
rect 1354 144 1355 148
rect 1359 144 1364 148
rect 1392 144 1393 148
rect 1397 144 1402 148
rect 1436 144 1437 148
rect 1441 144 1446 148
rect 1474 144 1475 148
rect 1479 144 1484 148
rect 1520 146 1521 150
rect 1525 146 1530 150
rect 286 85 295 143
rect 301 133 344 140
rect 378 133 385 143
rect 827 133 831 141
rect 855 133 859 141
rect 882 133 886 141
rect 921 133 925 141
rect 949 133 953 141
rect 976 133 980 141
rect 1016 134 1020 142
rect 1044 134 1048 142
rect 1071 134 1075 142
rect 1107 134 1111 142
rect 1360 138 1364 144
rect 1398 138 1402 144
rect 1442 138 1446 144
rect 1480 138 1484 144
rect 1526 140 1530 146
rect 1803 141 1807 146
rect 312 118 316 133
rect 372 129 399 133
rect 395 126 399 129
rect 286 81 313 85
rect 320 84 324 98
rect 361 87 365 106
rect 320 80 347 84
rect 320 78 324 80
rect 312 63 316 68
rect 301 56 337 63
rect 342 42 347 80
rect 361 75 365 81
rect 361 59 365 65
rect 369 75 373 106
rect 403 87 407 106
rect 389 82 396 86
rect 403 81 427 87
rect 403 75 407 81
rect 390 69 395 75
rect 369 58 373 65
rect 403 58 407 65
rect 369 54 407 58
rect 373 46 377 51
rect 342 34 383 42
rect 1792 134 1828 141
rect 1833 120 1838 158
rect 1852 153 1856 159
rect 1852 137 1856 143
rect 1860 153 1864 184
rect 1894 165 1898 184
rect 1880 160 1887 164
rect 1894 159 1918 165
rect 1894 153 1898 159
rect 1881 147 1886 153
rect 1860 136 1864 143
rect 1894 136 1898 143
rect 1860 132 1898 136
rect 1864 124 1868 129
rect 1833 112 1874 120
rect 1368 80 1372 98
rect 1406 80 1410 98
rect 1450 80 1454 98
rect 1488 80 1492 98
rect 1534 82 1538 100
rect 1851 88 1856 100
rect 1360 51 1364 60
rect 1398 51 1402 60
rect 1442 51 1446 60
rect 1480 51 1484 60
rect 1526 53 1530 62
rect 1360 47 1380 51
rect 1391 47 1422 51
rect 1434 47 1462 51
rect 1472 47 1489 51
rect 1509 49 1535 53
rect 835 27 839 33
rect 863 27 867 33
rect 890 27 894 33
rect 929 27 933 33
rect 957 27 961 33
rect 984 27 988 33
rect 1024 28 1028 34
rect 1052 28 1056 34
rect 1079 28 1083 34
rect 1115 28 1119 34
rect 360 10 365 22
rect 1840 5 1847 14
rect 43 -3 117 2
rect 43 -130 49 -3
rect 66 -13 99 -6
rect 113 -8 117 -3
rect 1874 -4 1881 12
rect 1782 -8 1881 -4
rect 77 -28 81 -13
rect 113 -15 142 -8
rect 55 -61 62 -58
rect 55 -65 78 -61
rect 85 -62 89 -48
rect 113 -61 120 -15
rect 112 -62 120 -61
rect 55 -112 60 -65
rect 85 -66 120 -62
rect 141 -64 145 -45
rect 85 -68 89 -66
rect 124 -70 145 -64
rect 141 -77 145 -70
rect 77 -83 81 -78
rect 66 -90 102 -83
rect 149 -63 153 -45
rect 149 -69 184 -63
rect 149 -77 153 -69
rect 116 -99 142 -92
rect 116 -112 123 -99
rect 55 -118 123 -112
rect 127 -108 135 -104
rect 127 -122 130 -108
rect 178 -112 184 -69
rect 1782 -66 1791 -8
rect 1797 -18 1840 -11
rect 1874 -18 1881 -8
rect 1808 -33 1812 -18
rect 1868 -22 1895 -18
rect 1891 -25 1895 -22
rect 1782 -70 1809 -66
rect 1816 -67 1820 -53
rect 1857 -64 1861 -45
rect 1816 -71 1843 -67
rect 1816 -73 1820 -71
rect 1808 -88 1812 -83
rect 1797 -95 1833 -88
rect 124 -126 130 -122
rect 140 -118 184 -112
rect 1838 -109 1843 -71
rect 1857 -76 1861 -70
rect 1857 -92 1861 -86
rect 1865 -76 1869 -45
rect 1899 -64 1903 -45
rect 1885 -69 1892 -65
rect 1899 -70 1923 -64
rect 1899 -76 1903 -70
rect 1886 -82 1891 -76
rect 1865 -93 1869 -86
rect 1899 -93 1903 -86
rect 1865 -97 1903 -93
rect 1869 -105 1873 -100
rect 1838 -117 1879 -109
rect 124 -130 127 -126
rect 140 -129 144 -118
rect 43 -134 127 -130
rect 132 -152 136 -139
rect 1856 -141 1861 -129
rect 120 -157 156 -152
rect 357 -177 364 -168
rect 391 -186 398 -170
rect 299 -190 398 -186
rect 299 -248 308 -190
rect 314 -200 357 -193
rect 391 -200 398 -190
rect 1840 -186 1847 -177
rect 1874 -195 1881 -179
rect 1782 -199 1881 -195
rect 325 -215 329 -200
rect 385 -204 412 -200
rect 408 -207 412 -204
rect 299 -252 326 -248
rect 333 -249 337 -235
rect 374 -246 378 -227
rect 333 -253 360 -249
rect 333 -255 337 -253
rect 325 -270 329 -265
rect 314 -277 350 -270
rect 355 -291 360 -253
rect 374 -258 378 -252
rect 374 -274 378 -268
rect 382 -258 386 -227
rect 416 -246 420 -227
rect 402 -251 409 -247
rect 416 -252 440 -246
rect 416 -258 420 -252
rect 403 -264 408 -258
rect 1782 -257 1791 -199
rect 1797 -209 1840 -202
rect 1874 -209 1881 -199
rect 1808 -224 1812 -209
rect 1868 -213 1895 -209
rect 1891 -216 1895 -213
rect 1782 -261 1809 -257
rect 1816 -258 1820 -244
rect 1857 -255 1861 -236
rect 1816 -262 1843 -258
rect 1816 -264 1820 -262
rect 382 -275 386 -268
rect 416 -275 420 -268
rect 382 -279 420 -275
rect 1808 -279 1812 -274
rect 386 -287 390 -282
rect 1797 -286 1833 -279
rect 355 -299 396 -291
rect 1838 -300 1843 -262
rect 1857 -267 1861 -261
rect 1857 -283 1861 -277
rect 1865 -267 1869 -236
rect 1899 -255 1903 -236
rect 1885 -260 1892 -256
rect 1899 -261 1923 -255
rect 1899 -267 1903 -261
rect 1886 -273 1891 -267
rect 1865 -284 1869 -277
rect 1899 -284 1903 -277
rect 1865 -288 1903 -284
rect 1869 -296 1873 -291
rect 1838 -308 1879 -300
rect 373 -323 378 -311
rect 1856 -332 1861 -320
rect 48 -377 122 -372
rect 48 -504 54 -377
rect 71 -387 104 -380
rect 118 -382 122 -377
rect 82 -402 86 -387
rect 118 -389 147 -382
rect 60 -435 67 -432
rect 60 -439 83 -435
rect 90 -436 94 -422
rect 118 -435 125 -389
rect 117 -436 125 -435
rect 60 -486 65 -439
rect 90 -440 125 -436
rect 146 -438 150 -419
rect 90 -442 94 -440
rect 129 -444 150 -438
rect 146 -451 150 -444
rect 82 -457 86 -452
rect 71 -464 107 -457
rect 154 -437 158 -419
rect 154 -443 189 -437
rect 154 -451 158 -443
rect 121 -473 147 -466
rect 121 -486 128 -473
rect 60 -492 128 -486
rect 132 -482 140 -478
rect 132 -496 135 -482
rect 183 -486 189 -443
rect 129 -500 135 -496
rect 145 -492 189 -486
rect 129 -504 132 -500
rect 145 -503 149 -492
rect 48 -508 132 -504
rect 137 -526 141 -513
rect 125 -531 161 -526
<< m2contact >>
rect 352 665 359 671
rect 352 648 359 655
rect 368 596 374 602
rect 368 569 373 574
rect 392 596 397 602
rect 391 584 398 590
rect 385 561 390 566
rect 391 549 398 557
rect 368 537 373 543
rect 1820 438 1827 444
rect 349 371 356 377
rect 349 354 356 361
rect 1820 421 1827 428
rect 365 302 371 308
rect 365 275 370 280
rect 1836 369 1842 375
rect 1836 342 1841 347
rect 1860 369 1865 375
rect 1859 357 1866 363
rect 1853 334 1858 339
rect 1859 322 1866 330
rect 389 302 394 308
rect 1836 310 1841 316
rect 388 290 395 296
rect 382 267 387 272
rect 388 255 395 263
rect 365 243 370 249
rect 1835 228 1842 234
rect 1835 211 1842 218
rect 344 150 351 156
rect 1851 159 1857 165
rect 344 133 351 140
rect 360 81 366 87
rect 360 54 365 59
rect 384 81 389 87
rect 383 69 390 75
rect 377 46 382 51
rect 383 34 390 42
rect 1851 132 1856 137
rect 1875 159 1880 165
rect 1874 147 1881 153
rect 1868 124 1873 129
rect 1874 112 1881 120
rect 1851 100 1856 106
rect 360 22 365 28
rect 1840 -1 1847 5
rect 1840 -18 1847 -11
rect 1856 -70 1862 -64
rect 1856 -97 1861 -92
rect 1880 -70 1885 -64
rect 1879 -82 1886 -76
rect 1873 -105 1878 -100
rect 1879 -117 1886 -109
rect 1856 -129 1861 -123
rect 357 -183 364 -177
rect 357 -200 364 -193
rect 1840 -192 1847 -186
rect 373 -252 379 -246
rect 373 -279 378 -274
rect 397 -252 402 -246
rect 396 -264 403 -258
rect 1840 -209 1847 -202
rect 1856 -261 1862 -255
rect 390 -287 395 -282
rect 396 -299 403 -291
rect 1856 -288 1861 -283
rect 1880 -261 1885 -255
rect 1879 -273 1886 -267
rect 1873 -296 1878 -291
rect 373 -311 378 -305
rect 1879 -308 1886 -300
rect 1856 -320 1861 -314
<< pm12contact >>
rect 890 296 896 302
rect 940 297 946 303
rect 990 297 996 303
rect 1037 297 1043 303
rect 1360 83 1365 88
rect 1398 83 1403 88
rect 1442 83 1447 88
rect 1480 83 1485 88
rect 1526 85 1531 90
rect 827 21 832 26
rect 855 21 860 26
rect 882 21 887 26
rect 921 21 926 26
rect 949 21 954 26
rect 976 21 981 26
rect 1016 22 1021 27
rect 1044 22 1049 27
rect 1071 22 1076 27
rect 1107 22 1112 27
<< metal2 >>
rect 352 655 359 665
rect 374 597 392 601
rect 368 543 373 569
rect 391 566 398 584
rect 390 561 398 566
rect 391 557 398 561
rect 1820 428 1827 438
rect 349 361 356 371
rect 1842 370 1860 374
rect 1836 316 1841 342
rect 1859 339 1866 357
rect 1858 334 1866 339
rect 1859 330 1866 334
rect 371 303 389 307
rect 880 296 890 302
rect 930 297 940 303
rect 980 297 990 303
rect 1027 297 1037 303
rect 365 249 370 275
rect 388 272 395 290
rect 387 267 395 272
rect 388 263 395 267
rect 1835 218 1842 228
rect 1857 160 1875 164
rect 344 140 351 150
rect 1851 106 1856 132
rect 1874 129 1881 147
rect 1873 124 1881 129
rect 1874 120 1881 124
rect 366 82 384 86
rect 1357 83 1360 88
rect 1395 83 1398 88
rect 1439 83 1442 88
rect 1477 83 1480 88
rect 1523 85 1526 90
rect 360 28 365 54
rect 383 51 390 69
rect 382 46 390 51
rect 383 42 390 46
rect 823 21 827 26
rect 851 21 855 26
rect 878 21 882 26
rect 917 21 921 26
rect 945 21 949 26
rect 972 21 976 26
rect 1012 22 1016 27
rect 1040 22 1044 27
rect 1067 22 1071 27
rect 1103 22 1107 27
rect 1840 -11 1847 -1
rect 1862 -69 1880 -65
rect 1856 -123 1861 -97
rect 1879 -100 1886 -82
rect 1878 -105 1886 -100
rect 1879 -109 1886 -105
rect 357 -193 364 -183
rect 1840 -202 1847 -192
rect 379 -251 397 -247
rect 1862 -260 1880 -256
rect 373 -305 378 -279
rect 396 -282 403 -264
rect 395 -287 403 -282
rect 396 -291 403 -287
rect 1856 -314 1861 -288
rect 1879 -291 1886 -273
rect 1878 -296 1886 -291
rect 1879 -300 1886 -296
<< labels >>
rlabel metal1 827 137 831 141 1 pdr1
rlabel metal2 823 21 827 26 2 prop_1
rlabel metal1 835 27 839 32 1 prop1_car0
rlabel metal1 855 136 859 141 1 prop1_car0
rlabel metal2 851 21 855 26 1 carry_0
rlabel metal1 863 27 867 32 1 clock_car0
rlabel metal1 882 136 886 141 1 clock_car0
rlabel metal2 878 21 882 26 1 clock_in
rlabel metal1 890 27 894 32 1 gnd!
rlabel metal1 921 136 925 141 1 pdr2
rlabel metal2 917 21 921 26 1 prop_2
rlabel metal1 929 27 933 32 1 pdr1
rlabel metal1 949 136 953 141 1 pdr1
rlabel metal2 945 21 949 26 1 gen_1
rlabel metal1 957 27 961 32 1 clock_car0
rlabel metal1 976 136 980 141 1 pdr3
rlabel metal2 972 21 976 26 1 prop_3
rlabel metal1 984 27 988 32 1 pdr2
rlabel metal1 1016 137 1020 142 1 pdr2
rlabel metal2 1012 22 1016 27 1 gen_2
rlabel metal1 1024 28 1028 33 1 clock_car0
rlabel metal1 1044 137 1048 142 1 pdr4
rlabel metal2 1040 22 1044 27 1 prop_4
rlabel metal1 1052 28 1056 33 1 pdr3
rlabel metal1 1071 137 1075 142 1 pdr3
rlabel metal2 1067 22 1071 27 1 gen_3
rlabel metal1 1079 28 1083 33 1 clock_car0
rlabel metal1 1107 137 1111 142 1 pdr4
rlabel metal2 1103 22 1107 27 1 gen_4
rlabel metal1 1115 28 1119 33 7 clock_car0
rlabel metal1 891 384 895 389 5 vdd!
rlabel metal1 941 385 945 390 5 vdd!
rlabel metal1 991 385 995 390 5 vdd!
rlabel metal1 1038 385 1042 390 5 vdd!
rlabel metal2 880 296 886 302 2 clock_in
rlabel metal2 930 297 936 303 1 clock_in
rlabel metal2 980 297 986 303 1 clock_in
rlabel metal2 1027 297 1032 303 1 clock_in
rlabel metal1 899 305 903 310 1 pdr1
rlabel metal1 949 306 953 310 1 pdr2
rlabel metal1 999 306 1003 310 1 pdr3
rlabel metal1 1046 306 1050 310 1 pdr4
rlabel metal1 1485 47 1489 51 1 gnd!
rlabel metal1 1481 151 1486 155 5 vdd!
rlabel metal2 1357 83 1360 88 1 pdr1
rlabel metal2 1395 83 1398 88 1 pdr2
rlabel metal2 1439 83 1442 88 1 pdr3
rlabel metal2 1477 83 1480 88 1 pdr4
rlabel metal1 1368 83 1372 88 1 c1
rlabel metal1 1406 83 1410 88 1 c2
rlabel metal1 1450 83 1454 88 1 c3
rlabel metal1 1488 83 1492 88 1 c4
rlabel metal1 1531 49 1535 53 1 gnd!
rlabel metal1 1527 153 1532 157 5 vdd!
rlabel metal2 1523 85 1526 90 1 clk_org
rlabel metal1 1534 85 1538 90 1 clock_in
rlabel metal1 1360 151 1364 155 5 vdd!
rlabel metal1 1398 151 1402 155 5 vdd!
rlabel metal1 1442 151 1446 155 5 vdd!
rlabel metal1 1446 47 1450 51 1 gnd!
rlabel metal1 1409 47 1413 51 1 gnd!
rlabel metal1 1369 47 1373 51 1 gnd!
rlabel metal2 1862 333 1862 333 1 bbar
rlabel metal1 1797 425 1797 425 1 vdd
rlabel metal1 1798 345 1798 345 1 gnd
rlabel metal1 1823 449 1823 449 5 vdd
rlabel metal1 1797 347 1797 347 1 gnd
rlabel metal1 1796 425 1796 425 5 vdd
rlabel metal1 1779 371 1779 371 1 invi
rlabel metal1 1815 370 1815 370 1 invo
rlabel metal2 1877 123 1877 123 1 bbar
rlabel metal1 1812 215 1812 215 1 vdd
rlabel metal1 1813 135 1813 135 1 gnd
rlabel metal1 1838 239 1838 239 5 vdd
rlabel metal1 1812 137 1812 137 1 gnd
rlabel metal1 1811 215 1811 215 5 vdd
rlabel metal1 1794 161 1794 161 1 invi
rlabel metal1 1830 160 1830 160 1 invo
rlabel metal2 1882 -106 1882 -106 1 bbar
rlabel metal1 1817 -14 1817 -14 1 vdd
rlabel metal1 1818 -94 1818 -94 1 gnd
rlabel metal1 1843 10 1843 10 5 vdd
rlabel metal1 1817 -92 1817 -92 1 gnd
rlabel metal1 1816 -14 1816 -14 5 vdd
rlabel metal1 1799 -68 1799 -68 1 invi
rlabel metal1 1835 -69 1835 -69 1 invo
rlabel metal2 1882 -297 1882 -297 1 bbar
rlabel metal1 1817 -205 1817 -205 1 vdd
rlabel metal1 1818 -285 1818 -285 1 gnd
rlabel metal1 1843 -181 1843 -181 5 vdd
rlabel metal1 1817 -283 1817 -283 1 gnd
rlabel metal1 1816 -205 1816 -205 5 vdd
rlabel metal1 1799 -259 1799 -259 1 invi
rlabel metal1 1835 -260 1835 -260 1 invo
rlabel metal2 394 560 394 560 1 bbar
rlabel metal1 329 652 329 652 1 vdd
rlabel metal1 330 572 330 572 1 gnd
rlabel metal1 355 676 355 676 5 vdd
rlabel metal1 329 574 329 574 1 gnd
rlabel metal1 328 652 328 652 5 vdd
rlabel metal1 311 598 311 598 1 invi
rlabel metal1 347 597 347 597 1 invo
rlabel metal2 386 45 386 45 1 bbar
rlabel metal1 321 137 321 137 1 vdd
rlabel metal1 322 57 322 57 1 gnd
rlabel metal1 347 161 347 161 5 vdd
rlabel metal1 321 59 321 59 1 gnd
rlabel metal1 320 137 320 137 5 vdd
rlabel metal1 303 83 303 83 1 invi
rlabel metal1 339 82 339 82 1 invo
rlabel metal2 399 -288 399 -288 1 bbar
rlabel metal1 334 -196 334 -196 1 vdd
rlabel metal1 335 -276 335 -276 1 gnd
rlabel metal1 360 -172 360 -172 5 vdd
rlabel metal1 334 -274 334 -274 1 gnd
rlabel metal1 333 -196 333 -196 5 vdd
rlabel metal1 316 -250 316 -250 1 invi
rlabel metal1 352 -251 352 -251 1 invo
rlabel metal2 391 266 391 266 1 bbar
rlabel metal1 326 358 326 358 1 vdd
rlabel metal1 327 278 327 278 1 gnd
rlabel metal1 352 382 352 382 5 vdd
rlabel metal1 326 280 326 280 1 gnd
rlabel metal1 325 358 325 358 5 vdd
rlabel metal1 308 304 308 304 1 invi
rlabel metal1 344 303 344 303 1 invo
rlabel metal1 378 155 385 163 1 q_b1
rlabel metal1 360 10 365 17 1 q_a1
rlabel metal1 420 82 427 87 1 prop_1
rlabel metal1 391 -177 398 -170 1 q_b2
rlabel metal1 373 -323 378 -316 1 q_a2
rlabel metal1 434 -252 440 -246 1 prop_2
rlabel metal1 383 376 390 384 1 q_b3
rlabel metal1 425 302 432 308 1 prop_3
rlabel metal1 365 231 370 238 1 q_a3
rlabel metal1 386 670 393 678 1 q_b4
rlabel metal1 368 525 373 532 1 q_a4
rlabel metal1 429 596 435 602 1 prop_4
rlabel metal1 1836 298 1841 305 1 prop_1
rlabel metal1 1897 369 1903 375 1 s1
rlabel metal1 1851 88 1856 96 1 prop_2
rlabel metal1 1911 159 1918 165 1 s2
rlabel metal1 1854 442 1861 451 1 carry_0
rlabel metal1 1869 233 1876 241 1 c1
rlabel metal1 1874 4 1881 12 1 c2
rlabel metal1 1856 -141 1861 -133 1 prop_3
rlabel metal1 1916 -70 1923 -64 7 s3
rlabel metal1 1874 -186 1881 -179 1 c3
rlabel metal1 1856 -332 1861 -325 1 prop_4
rlabel metal1 1917 -261 1923 -255 7 s4
rlabel metal1 150 504 150 504 1 invo
rlabel metal1 114 505 114 505 1 invi
rlabel metal1 131 559 131 559 5 vdd
rlabel metal1 132 481 132 481 1 gnd
rlabel metal1 105 222 105 222 1 gnd
rlabel metal1 104 300 104 300 5 vdd
rlabel metal1 87 246 87 246 1 invi
rlabel metal1 123 245 123 245 1 invo
rlabel metal1 104 -64 104 -64 1 invo
rlabel metal1 68 -63 68 -63 1 invi
rlabel metal1 85 -9 85 -9 5 vdd
rlabel metal1 86 -87 86 -87 1 gnd
rlabel metal1 109 -438 109 -438 1 invo
rlabel metal1 73 -437 73 -437 1 invi
rlabel metal1 90 -383 90 -383 5 vdd
rlabel metal1 91 -461 91 -461 1 gnd
rlabel metal1 170 498 176 504 1 q_a1
rlabel metal1 162 469 170 475 1 q_b1
rlabel metal1 224 491 230 496 1 gen_1
rlabel metal1 143 239 152 245 1 q_a2
rlabel metal1 135 210 144 216 1 q_b2
rlabel metal1 193 240 202 246 1 gen_2
rlabel metal1 124 -70 133 -64 1 q_a3
rlabel metal1 116 -99 125 -93 1 q_b3
rlabel metal1 175 -69 184 -63 1 gen_3
rlabel metal1 129 -444 138 -438 1 q_a4
rlabel metal1 121 -473 130 -467 1 q_b4
rlabel metal1 179 -443 188 -437 1 gen_4
<< end >>
