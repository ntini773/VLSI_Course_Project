magic
tech scmos
timestamp 1732012043
<< nwell >>
rect 13 -87 45 -50
rect 51 -87 77 -50
rect 95 -87 121 -50
rect 140 -87 166 -50
<< ntransistor >>
rect 20 -113 22 -103
rect 56 -113 58 -103
rect 64 -113 66 -103
rect 100 -113 102 -103
rect 108 -113 110 -103
rect 151 -113 153 -103
<< ptransistor >>
rect 24 -81 26 -56
rect 32 -81 34 -56
rect 62 -81 64 -56
rect 106 -81 108 -56
rect 151 -81 153 -56
<< ndiffusion >>
rect 19 -113 20 -103
rect 22 -113 23 -103
rect 55 -113 56 -103
rect 58 -113 59 -103
rect 63 -113 64 -103
rect 66 -113 67 -103
rect 99 -113 100 -103
rect 102 -113 103 -103
rect 107 -113 108 -103
rect 110 -113 111 -103
rect 150 -113 151 -103
rect 153 -113 154 -103
<< pdiffusion >>
rect 23 -81 24 -56
rect 26 -81 27 -56
rect 31 -81 32 -56
rect 34 -81 35 -56
rect 61 -81 62 -56
rect 64 -81 65 -56
rect 105 -81 106 -56
rect 108 -81 109 -56
rect 150 -81 151 -56
rect 153 -81 154 -56
<< ndcontact >>
rect 15 -113 19 -103
rect 23 -113 27 -103
rect 51 -113 55 -103
rect 59 -113 63 -103
rect 67 -113 71 -103
rect 95 -113 99 -103
rect 103 -113 107 -103
rect 111 -113 115 -103
rect 146 -113 150 -103
rect 154 -113 158 -103
<< pdcontact >>
rect 19 -81 23 -56
rect 27 -81 31 -56
rect 35 -81 39 -56
rect 57 -81 61 -56
rect 65 -81 69 -56
rect 101 -81 105 -56
rect 109 -81 113 -56
rect 146 -81 150 -56
rect 154 -81 158 -56
<< polysilicon >>
rect 24 -56 26 -53
rect 32 -56 34 -53
rect 62 -56 64 -53
rect 106 -56 108 -53
rect 151 -56 153 -53
rect 24 -88 26 -81
rect 19 -92 26 -88
rect 20 -103 22 -92
rect 32 -100 34 -81
rect 62 -89 64 -81
rect 106 -89 108 -81
rect 56 -91 64 -89
rect 100 -91 108 -89
rect 56 -103 58 -91
rect 64 -103 66 -94
rect 100 -103 102 -91
rect 108 -103 110 -94
rect 151 -103 153 -81
rect 20 -116 22 -113
rect 56 -116 58 -113
rect 64 -116 66 -113
rect 100 -116 102 -113
rect 108 -116 110 -113
rect 151 -116 153 -113
<< polycontact >>
rect 15 -92 19 -88
rect 28 -100 32 -96
rect 51 -100 56 -95
rect 66 -100 71 -96
rect 95 -100 100 -95
rect 147 -95 151 -90
rect 110 -100 115 -96
<< metal1 >>
rect 13 -50 166 -46
rect 19 -56 23 -50
rect 57 -56 61 -50
rect 101 -56 105 -50
rect 146 -56 150 -50
rect 69 -81 82 -56
rect 113 -81 126 -56
rect 8 -92 15 -88
rect 35 -89 39 -81
rect 35 -95 43 -89
rect 79 -90 82 -81
rect 123 -90 126 -81
rect 79 -95 87 -90
rect 123 -95 147 -90
rect 154 -91 158 -81
rect 25 -100 28 -96
rect 35 -103 39 -95
rect 47 -100 51 -95
rect 71 -100 75 -96
rect 79 -103 82 -95
rect 91 -100 95 -95
rect 115 -100 119 -96
rect 123 -103 126 -95
rect 154 -96 167 -91
rect 154 -103 158 -96
rect 27 -113 39 -103
rect 71 -113 82 -103
rect 115 -113 126 -103
rect 15 -118 19 -113
rect 51 -118 55 -113
rect 95 -118 99 -113
rect 146 -118 150 -113
rect 14 -122 158 -118
<< labels >>
rlabel metal1 23 -120 26 -119 1 gnd
rlabel metal1 40 -92 41 -91 1 x
rlabel metal1 72 -99 74 -97 7 x
rlabel metal1 84 -93 85 -92 7 y
rlabel metal1 92 -99 93 -97 1 y
rlabel metal1 128 -93 129 -92 1 qb
rlabel metal1 26 -98 26 -98 1 clk_org
rlabel metal1 49 -97 49 -97 1 clk_org
rlabel metal1 117 -97 117 -97 1 clk_org
rlabel metal1 34 -48 34 -48 5 vdd
<< end >>
