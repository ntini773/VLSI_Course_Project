magic
tech scmos
timestamp 1731618937
<< nwell >>
rect -17 -22 16 25
<< ntransistor >>
rect -1 -40 1 -30
<< ptransistor >>
rect -1 -10 1 10
<< ndiffusion >>
rect -2 -40 -1 -30
rect 1 -40 2 -30
<< pdiffusion >>
rect -2 -10 -1 10
rect 1 -10 2 10
<< ndcontact >>
rect -6 -40 -2 -30
rect 2 -40 6 -30
<< pdcontact >>
rect -6 -10 -2 10
rect 2 -10 6 10
<< polysilicon >>
rect -1 10 1 19
rect -1 -30 1 -10
rect -1 -43 1 -40
<< polycontact >>
rect -5 -27 -1 -23
<< metal1 >>
rect -17 25 16 32
rect -6 10 -2 25
rect -23 -27 -5 -23
rect 2 -24 6 -10
rect 2 -28 29 -24
rect 2 -30 6 -28
rect -6 -45 -2 -40
rect -17 -52 19 -45
<< labels >>
rlabel metal1 3 -49 3 -49 1 gnd
rlabel metal1 2 29 2 29 5 vdd
rlabel metal1 -15 -25 -15 -25 1 invi
rlabel metal1 21 -26 21 -26 1 invo
<< end >>
