magic
tech scmos
timestamp 1732103492
<< nwell >>
rect 2033 928 2085 952
rect 2200 885 2252 909
rect 2382 878 2434 902
rect 2668 754 2692 806
rect 2539 723 2601 747
rect 1995 661 2057 685
rect 2169 684 2231 708
rect 2343 688 2405 712
rect 2067 369 2119 393
rect 1876 340 1913 366
rect 1876 295 1913 321
rect 1876 251 1913 277
rect 1876 213 1913 245
<< ntransistor >>
rect 2097 939 2117 941
rect 2264 896 2284 898
rect 2446 889 2466 891
rect 2679 722 2681 742
rect 2521 649 2621 651
rect 2333 641 2433 643
rect 2152 631 2252 633
rect 1984 623 2084 625
rect 2523 540 2623 542
rect 2331 530 2431 532
rect 2151 520 2251 522
rect 1936 412 1938 512
rect 1983 509 2083 511
rect 2016 411 2116 413
rect 2131 380 2151 382
rect 1929 351 1939 353
rect 1929 308 1939 310
rect 1929 300 1939 302
rect 1929 264 1939 266
rect 1929 256 1939 258
rect 1929 220 1939 222
<< ptransistor >>
rect 2039 939 2079 941
rect 2206 896 2246 898
rect 2388 889 2428 891
rect 2679 760 2681 800
rect 2545 734 2595 736
rect 2349 699 2399 701
rect 2175 695 2225 697
rect 2001 672 2051 674
rect 2073 380 2113 382
rect 1882 351 1907 353
rect 1882 306 1907 308
rect 1882 262 1907 264
rect 1882 232 1907 234
rect 1882 224 1907 226
<< ndiffusion >>
rect 2097 941 2117 942
rect 2097 938 2117 939
rect 2264 898 2284 899
rect 2264 895 2284 896
rect 2446 891 2466 892
rect 2446 888 2466 889
rect 2678 722 2679 742
rect 2681 722 2682 742
rect 2521 651 2621 652
rect 2521 648 2621 649
rect 2333 643 2433 644
rect 2333 640 2433 641
rect 2152 633 2252 634
rect 2152 630 2252 631
rect 1984 625 2084 626
rect 1984 622 2084 623
rect 2523 542 2623 543
rect 2523 539 2623 540
rect 2331 532 2431 533
rect 2331 529 2431 530
rect 2151 522 2251 523
rect 2151 519 2251 520
rect 1935 412 1936 512
rect 1938 412 1939 512
rect 1983 511 2083 512
rect 1983 508 2083 509
rect 2016 413 2116 414
rect 2016 410 2116 411
rect 2131 382 2151 383
rect 2131 379 2151 380
rect 1929 353 1939 354
rect 1929 350 1939 351
rect 1929 310 1939 311
rect 1929 307 1939 308
rect 1929 302 1939 303
rect 1929 299 1939 300
rect 1929 266 1939 267
rect 1929 263 1939 264
rect 1929 258 1939 259
rect 1929 255 1939 256
rect 1929 222 1939 223
rect 1929 219 1939 220
<< pdiffusion >>
rect 2039 941 2079 942
rect 2039 938 2079 939
rect 2206 898 2246 899
rect 2206 895 2246 896
rect 2388 891 2428 892
rect 2388 888 2428 889
rect 2678 760 2679 800
rect 2681 760 2682 800
rect 2545 736 2595 737
rect 2545 733 2595 734
rect 2175 697 2225 698
rect 2349 701 2399 702
rect 2349 698 2399 699
rect 2175 694 2225 695
rect 2001 674 2051 675
rect 2001 671 2051 672
rect 2073 382 2113 383
rect 2073 379 2113 380
rect 1882 353 1907 354
rect 1882 350 1907 351
rect 1882 308 1907 309
rect 1882 305 1907 306
rect 1882 264 1907 265
rect 1882 261 1907 262
rect 1882 234 1907 235
rect 1882 231 1907 232
rect 1882 226 1907 227
rect 1882 223 1907 224
<< ndcontact >>
rect 2097 942 2117 946
rect 2097 934 2117 938
rect 2264 899 2284 903
rect 2264 891 2284 895
rect 2446 892 2466 896
rect 2446 884 2466 888
rect 2674 722 2678 742
rect 2682 722 2686 742
rect 2521 652 2621 656
rect 2333 644 2433 648
rect 2521 644 2621 648
rect 2152 634 2252 638
rect 2333 636 2433 640
rect 1984 626 2084 630
rect 2152 626 2252 630
rect 1984 618 2084 622
rect 2523 543 2623 547
rect 2331 533 2431 537
rect 2523 535 2623 539
rect 2151 523 2251 527
rect 2331 525 2431 529
rect 1931 412 1935 512
rect 1939 412 1943 512
rect 1983 512 2083 516
rect 2151 515 2251 519
rect 1983 504 2083 508
rect 2016 414 2116 418
rect 2016 406 2116 410
rect 2131 383 2151 387
rect 2131 375 2151 379
rect 1929 354 1939 358
rect 1929 346 1939 350
rect 1929 311 1939 315
rect 1929 303 1939 307
rect 1929 295 1939 299
rect 1929 267 1939 271
rect 1929 259 1939 263
rect 1929 251 1939 255
rect 1929 223 1939 227
rect 1929 215 1939 219
<< pdcontact >>
rect 2039 942 2079 946
rect 2039 934 2079 938
rect 2206 899 2246 903
rect 2206 891 2246 895
rect 2388 892 2428 896
rect 2388 884 2428 888
rect 2674 760 2678 800
rect 2682 760 2686 800
rect 2545 737 2595 741
rect 2545 729 2595 733
rect 2175 698 2225 702
rect 2349 702 2399 706
rect 2349 694 2399 698
rect 2175 690 2225 694
rect 2001 675 2051 679
rect 2001 667 2051 671
rect 2073 383 2113 387
rect 2073 375 2113 379
rect 1882 354 1907 358
rect 1882 346 1907 350
rect 1882 309 1907 313
rect 1882 301 1907 305
rect 1882 265 1907 269
rect 1882 257 1907 261
rect 1882 235 1907 239
rect 1882 227 1907 231
rect 1882 219 1907 223
<< nsubstratencontact >>
rect 2029 929 2033 933
rect 2196 886 2200 890
rect 2378 879 2382 883
rect 2669 806 2673 810
rect 2534 742 2539 746
rect 2338 707 2343 711
rect 2164 703 2169 707
rect 1990 680 1995 684
rect 2063 370 2067 374
<< polysilicon >>
rect 2036 939 2039 941
rect 2079 939 2097 941
rect 2117 939 2121 941
rect 2203 896 2206 898
rect 2246 896 2264 898
rect 2284 896 2288 898
rect 2385 889 2388 891
rect 2428 889 2446 891
rect 2466 889 2470 891
rect 2679 800 2681 803
rect 2679 742 2681 760
rect 2542 734 2545 736
rect 2595 734 2618 736
rect 2679 718 2681 722
rect 2346 699 2349 701
rect 2399 699 2422 701
rect 2172 695 2175 697
rect 2225 695 2248 697
rect 1998 672 2001 674
rect 2051 672 2074 674
rect 2509 649 2521 651
rect 2621 649 2624 651
rect 2321 641 2333 643
rect 2433 641 2436 643
rect 2140 631 2152 633
rect 2252 631 2255 633
rect 1972 623 1984 625
rect 2084 623 2087 625
rect 2511 540 2523 542
rect 2623 540 2626 542
rect 2319 530 2331 532
rect 2431 530 2434 532
rect 2139 520 2151 522
rect 2251 520 2254 522
rect 1936 512 1938 515
rect 1971 509 1983 511
rect 2083 509 2086 511
rect 1936 400 1938 412
rect 2013 411 2016 413
rect 2116 411 2128 413
rect 2070 380 2073 382
rect 2113 380 2131 382
rect 2151 380 2155 382
rect 1879 351 1882 353
rect 1907 351 1929 353
rect 1939 351 1942 353
rect 1920 308 1929 310
rect 1939 308 1942 310
rect 1879 306 1882 308
rect 1907 306 1917 308
rect 1915 302 1917 306
rect 1915 300 1929 302
rect 1939 300 1942 302
rect 1920 264 1929 266
rect 1939 264 1942 266
rect 1879 262 1882 264
rect 1907 262 1917 264
rect 1915 258 1917 262
rect 1915 256 1929 258
rect 1939 256 1942 258
rect 1879 232 1882 234
rect 1907 232 1926 234
rect 1879 224 1882 226
rect 1907 224 1918 226
rect 1914 222 1918 224
rect 1914 220 1929 222
rect 1939 220 1942 222
rect 1914 219 1918 220
<< polycontact >>
rect 2674 745 2679 750
rect 1916 347 1921 351
rect 1922 310 1926 314
rect 1921 295 1926 300
rect 1922 266 1926 270
rect 1921 251 1926 256
rect 1914 239 1918 243
rect 1922 228 1926 232
rect 1914 215 1918 219
<< metal1 >>
rect 1898 413 1901 1050
rect 2022 938 2026 954
rect 2087 946 2090 1050
rect 2079 942 2097 946
rect 2022 934 2039 938
rect 2126 938 2130 954
rect 2117 934 2130 938
rect 2029 933 2033 934
rect 2029 928 2033 929
rect 1990 684 1995 685
rect 1990 679 1995 680
rect 1981 675 2001 679
rect 1990 661 1995 675
rect 2089 671 2093 902
rect 2189 895 2193 915
rect 2256 903 2259 921
rect 2246 899 2264 903
rect 2189 891 2206 895
rect 2293 895 2297 915
rect 2284 891 2297 895
rect 2189 884 2193 891
rect 2196 890 2200 891
rect 2196 885 2200 886
rect 2293 884 2297 891
rect 2371 888 2375 904
rect 2439 896 2442 921
rect 2428 892 2446 896
rect 2371 884 2388 888
rect 2475 888 2479 904
rect 2466 884 2479 888
rect 2371 876 2375 884
rect 2378 883 2382 884
rect 2378 878 2382 879
rect 2475 876 2479 884
rect 2256 852 2261 858
rect 2164 707 2169 708
rect 2164 702 2169 703
rect 2155 698 2175 702
rect 2164 684 2169 698
rect 2257 694 2261 852
rect 2438 841 2443 845
rect 2439 826 2442 841
rect 2338 711 2343 712
rect 2338 706 2343 707
rect 2329 702 2349 706
rect 2225 690 2261 694
rect 2051 667 2093 671
rect 2089 630 2093 667
rect 2257 640 2261 690
rect 2338 688 2343 702
rect 2438 698 2442 826
rect 2666 813 2687 817
rect 2674 810 2678 813
rect 2668 806 2669 810
rect 2673 806 2678 810
rect 2674 800 2678 806
rect 2534 746 2539 747
rect 2628 745 2674 750
rect 2682 749 2686 760
rect 2682 745 2696 749
rect 2534 741 2539 742
rect 2525 737 2545 741
rect 2534 723 2539 737
rect 2628 733 2632 745
rect 2682 742 2686 745
rect 2595 729 2632 733
rect 2399 694 2442 698
rect 2438 648 2442 694
rect 2628 656 2632 729
rect 2674 713 2678 722
rect 2666 709 2683 713
rect 2621 652 2632 656
rect 2433 644 2521 648
rect 2256 638 2333 640
rect 2252 636 2333 638
rect 2252 634 2260 636
rect 2084 626 2152 630
rect 1882 408 1901 413
rect 1931 618 1984 622
rect 1931 512 1935 618
rect 2089 516 2093 626
rect 2256 527 2260 634
rect 2437 537 2441 644
rect 2628 547 2632 652
rect 2623 543 2632 547
rect 2431 533 2441 537
rect 2516 535 2523 539
rect 2251 523 2260 527
rect 2325 525 2331 529
rect 2083 512 2093 516
rect 2145 515 2151 519
rect 1977 504 1983 508
rect 1882 389 1887 408
rect 1898 405 1901 408
rect 1939 410 1943 412
rect 1978 499 1982 504
rect 2145 499 2149 515
rect 2325 499 2329 525
rect 2516 499 2520 535
rect 1978 495 2520 499
rect 1978 410 1982 495
rect 2116 414 2122 418
rect 1939 406 2016 410
rect 1882 384 1922 389
rect 1872 350 1876 366
rect 1917 358 1922 384
rect 2056 379 2060 388
rect 2113 385 2123 387
rect 2128 385 2131 387
rect 2113 383 2131 385
rect 2056 375 2073 379
rect 2160 379 2164 384
rect 2151 375 2164 379
rect 2056 365 2060 375
rect 2063 374 2067 375
rect 2063 369 2067 370
rect 2160 366 2164 375
rect 1907 354 1929 358
rect 1872 346 1882 350
rect 1944 350 1948 358
rect 1872 305 1876 346
rect 1916 326 1921 347
rect 1939 346 1948 350
rect 1882 323 1939 326
rect 1882 313 1907 323
rect 1922 314 1926 315
rect 1929 315 1939 323
rect 1872 301 1882 305
rect 1872 261 1876 301
rect 1944 299 1948 346
rect 1939 295 1948 299
rect 1921 291 1926 295
rect 1916 287 1926 291
rect 1916 282 1921 287
rect 1882 279 1939 282
rect 1882 269 1907 279
rect 1922 270 1926 271
rect 1929 271 1939 279
rect 1872 257 1882 261
rect 1872 223 1876 257
rect 1944 255 1948 295
rect 1939 251 1948 255
rect 1914 243 1918 244
rect 1921 248 1926 251
rect 1921 243 1923 248
rect 1907 235 1939 239
rect 1872 219 1882 223
rect 1922 219 1926 228
rect 1929 227 1939 235
rect 1944 219 1948 251
rect 1872 213 1876 219
rect 1914 208 1918 215
rect 1939 215 1948 219
rect 1944 214 1948 215
rect 1830 116 1839 120
<< m2contact >>
rect 2089 902 2094 908
rect 2256 858 2261 866
rect 2438 845 2443 851
rect 1898 400 1903 405
rect 2123 385 2128 390
rect 1921 315 1926 320
rect 1921 271 1926 276
rect 1913 244 1918 249
rect 1923 243 1928 248
rect 1921 214 1926 219
rect 1839 116 1844 122
<< pm12contact >>
rect 2089 934 2094 939
rect 2068 674 2074 680
rect 2256 891 2261 896
rect 2438 884 2443 889
rect 2242 697 2248 703
rect 2416 701 2422 707
rect 2612 736 2618 742
rect 2509 651 2514 656
rect 2321 643 2326 648
rect 2140 633 2145 638
rect 1972 625 1977 630
rect 2511 542 2516 547
rect 2319 532 2324 537
rect 2139 522 2144 527
rect 1971 511 1976 516
rect 2123 406 2128 411
rect 1931 400 1936 405
rect 2123 375 2128 380
<< metal2 >>
rect 1830 1017 1854 1022
rect 1830 887 1842 892
rect 1837 598 1842 887
rect 1849 613 1854 1017
rect 1972 638 1977 1050
rect 2089 908 2094 934
rect 2068 680 2074 684
rect 2140 648 2145 1050
rect 2256 866 2261 891
rect 2242 703 2248 707
rect 2321 657 2325 921
rect 2438 851 2443 884
rect 2493 832 2498 921
rect 2493 827 2514 832
rect 2493 826 2498 827
rect 2416 707 2422 711
rect 2509 669 2514 827
rect 2612 742 2618 746
rect 1962 633 1977 638
rect 1962 613 1967 633
rect 1972 630 1977 633
rect 2131 643 2145 648
rect 1849 608 1967 613
rect 2131 598 2136 643
rect 2140 638 2145 643
rect 2312 653 2325 657
rect 1837 593 2136 598
rect 2312 588 2316 653
rect 2321 652 2325 653
rect 2496 664 2514 669
rect 2321 648 2326 652
rect 1830 584 2316 588
rect 2496 578 2501 664
rect 2509 656 2514 664
rect 1830 573 2501 578
rect 1830 549 2516 554
rect 2511 547 2516 549
rect 1830 539 2324 544
rect 2319 537 2324 539
rect 1836 528 2144 534
rect 2139 527 2144 528
rect 1839 519 1976 524
rect 1839 122 1844 519
rect 1971 516 1976 519
rect 1903 400 1931 405
rect 2123 400 2128 406
rect 2123 390 2128 395
rect 2123 372 2128 375
rect 1950 320 1953 324
rect 1926 315 1953 320
rect 1865 271 1921 275
rect 1865 248 1869 271
rect 1865 244 1913 248
rect 1950 248 1953 315
rect 1928 244 1953 248
rect 1922 211 1926 214
rect 1950 211 1953 244
rect 1922 205 1953 211
rect 1922 193 1926 205
<< m3contact >>
rect 2068 684 2074 690
rect 2242 707 2248 713
rect 2416 711 2422 717
rect 2612 746 2618 752
rect 2123 395 2128 400
<< metal3 >>
rect 2068 777 2618 782
rect 2068 690 2074 777
rect 2242 713 2248 777
rect 2280 400 2285 777
rect 2416 717 2422 777
rect 2612 752 2618 777
rect 2128 395 2285 400
<< labels >>
rlabel metal1 2086 512 2091 516 3 pdr1
rlabel metal2 1971 516 1976 520 3 gen_1
rlabel metal1 1931 515 1935 520 1 prop1_car0
rlabel metal2 1927 400 1931 405 1 carry_0
rlabel metal1 1939 406 1943 411 1 clock_car0
rlabel metal1 2008 406 2013 410 7 clock_car0
rlabel metal2 2123 402 2128 406 7 clock_in
rlabel metal1 2117 414 2122 418 7 gnd!
rlabel metal1 1977 504 1982 508 3 clock_car0
rlabel metal1 2088 626 2092 630 3 pdr1
rlabel metal2 1972 630 1977 634 4 prop_1
rlabel metal1 1978 618 1983 622 3 prop1_car0
rlabel metal1 1981 675 1986 679 3 vdd!
rlabel m3contact 2068 684 2074 690 6 clock_in
rlabel metal1 2060 667 2065 671 7 pdr1
rlabel metal1 2145 515 2150 519 3 clock_car0
rlabel metal2 2139 527 2144 531 3 gen_2
rlabel metal1 2254 523 2259 527 3 pdr2
rlabel metal1 2255 634 2260 638 3 pdr2
rlabel metal2 2140 638 2145 642 3 prop_2
rlabel metal1 2146 626 2151 630 3 pdr1
rlabel metal1 2155 698 2160 702 3 vdd!
rlabel m3contact 2242 707 2248 713 7 clock_in
rlabel metal1 2235 690 2239 694 7 pdr2
rlabel metal1 2325 525 2330 529 3 clock_car0
rlabel metal2 2319 537 2324 541 3 gen_3
rlabel metal1 2434 533 2439 537 3 pdr3
rlabel metal1 2626 543 2631 547 3 pdr4
rlabel metal2 2511 547 2516 551 3 gen_4
rlabel metal1 2517 535 2522 539 1 clock_car0
rlabel metal1 2436 644 2441 648 3 pdr3
rlabel metal2 2321 648 2326 652 3 prop_3
rlabel metal1 2327 636 2332 640 3 pdr2
rlabel metal1 2624 652 2629 656 3 pdr4
rlabel metal2 2509 656 2514 660 3 prop_4
rlabel metal1 2515 644 2520 648 3 pdr3
rlabel metal1 2329 702 2334 706 3 vdd!
rlabel m3contact 2416 711 2422 717 7 clock_in
rlabel metal1 2409 694 2413 698 7 pdr3
rlabel metal1 2525 737 2530 741 3 vdd!
rlabel m3contact 2612 747 2618 752 7 clock_in
rlabel metal1 2605 729 2609 733 7 pdr4
rlabel metal1 2682 745 2686 750 1 c4
rlabel metal1 2675 813 2680 817 5 vdd!
rlabel metal1 2679 709 2683 713 1 gnd!
rlabel metal1 2160 380 2164 384 7 gnd!
rlabel metal1 2056 376 2060 381 3 vdd!
rlabel metal2 2123 372 2128 375 7 clk_org
rlabel metal1 2123 383 2128 387 7 clock_in
rlabel metal1 1945 223 1946 226 7 gnd
rlabel metal1 1873 229 1874 231 3 vdd
rlabel metal2 1925 210 1925 210 7 clk_org
rlabel metal1 1916 209 1916 209 7 cin
rlabel metal1 1920 366 1920 366 7 carry_0
rlabel metal2 2438 881 2443 884 7 pdr3
rlabel metal1 2438 892 2443 896 7 c3
rlabel metal1 2371 884 2375 888 3 vdd!
rlabel metal1 2475 888 2479 892 7 gnd!
rlabel metal1 2293 902 2297 906 7 gnd!
rlabel metal1 2189 891 2193 895 3 vdd!
rlabel metal1 2256 899 2261 903 7 c2
rlabel metal2 2256 888 2261 891 7 pdr2
rlabel metal2 2089 931 2094 934 7 pdr1
rlabel metal1 2089 942 2094 946 7 c1
rlabel metal1 2022 934 2026 938 3 vdd!
rlabel metal1 2126 943 2130 947 7 gnd!
<< end >>
