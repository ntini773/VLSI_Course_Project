magic
tech scmos
timestamp 1732061603
<< nwell >>
rect 4120 1202 4152 1226
rect 4115 1162 4152 1188
rect 3647 1108 3684 1140
rect 4115 1117 4152 1143
rect 4307 1141 4339 1165
rect 3647 1076 3684 1102
rect 4115 1073 4152 1099
rect 4302 1093 4339 1119
rect 4484 1117 4516 1141
rect 3548 1036 3585 1068
rect 3647 1032 3684 1058
rect 4115 1035 4152 1067
rect 4302 1048 4339 1074
rect 4479 1070 4516 1096
rect 3548 1004 3585 1030
rect 3647 987 3684 1013
rect 3908 1002 3940 1026
rect 4302 1004 4339 1030
rect 4479 1025 4516 1051
rect 3452 948 3489 980
rect 3548 960 3585 986
rect 3688 955 3712 979
rect 3727 969 3761 975
rect 3350 907 3387 939
rect 3452 916 3489 942
rect 3548 915 3585 941
rect 3727 939 3789 969
rect 3903 953 3940 979
rect 4070 948 4106 976
rect 4302 966 4339 998
rect 4479 981 4516 1007
rect 3755 933 3789 939
rect 4064 942 4106 948
rect 4479 943 4516 975
rect 3350 875 3387 901
rect 3688 900 3712 924
rect 3903 908 3940 934
rect 4064 914 4100 942
rect 4239 904 4275 932
rect 3452 872 3489 898
rect 3903 864 3940 890
rect 4060 875 4084 899
rect 4115 875 4139 899
rect 4233 898 4275 904
rect 4233 870 4269 898
rect 4422 874 4458 902
rect 4416 868 4458 874
rect 3246 810 3283 842
rect 3350 831 3387 857
rect 3452 827 3489 853
rect 3689 823 3713 847
rect 3728 837 3762 843
rect 3149 775 3186 807
rect 3246 778 3283 804
rect 3350 786 3387 812
rect 3728 807 3790 837
rect 3903 826 3940 858
rect 4229 831 4253 855
rect 4284 831 4308 855
rect 4416 840 4452 868
rect 3756 801 3790 807
rect 3149 743 3186 769
rect 3689 768 3713 792
rect 3246 734 3283 760
rect 3879 759 3915 787
rect 4033 785 4085 809
rect 4412 801 4436 825
rect 4467 801 4491 825
rect 3873 753 3915 759
rect 3047 702 3084 734
rect 3873 725 3909 753
rect 4200 742 4252 766
rect 4382 735 4434 759
rect 3149 699 3186 725
rect 2940 645 2977 677
rect 3047 670 3084 696
rect 3246 689 3283 715
rect 3149 654 3186 680
rect 3692 679 3716 703
rect 3731 693 3765 699
rect 3731 663 3793 693
rect 3869 686 3893 710
rect 3924 686 3948 710
rect 3759 657 3793 663
rect 2940 613 2977 639
rect 3047 626 3084 652
rect 3692 624 3716 648
rect 4668 611 4692 663
rect 4715 607 4747 644
rect 4753 607 4779 644
rect 4797 607 4823 644
rect 4842 607 4868 644
rect 2940 569 2977 595
rect 3047 581 3084 607
rect 4880 604 4904 636
rect 4539 580 4601 604
rect 3699 554 3723 578
rect 3738 568 3772 574
rect 2940 524 2977 550
rect 3738 538 3800 568
rect 3766 532 3800 538
rect 3699 499 3723 523
rect 3995 518 4057 542
rect 4169 541 4231 565
rect 4343 545 4405 569
rect 3721 321 3757 361
rect 3763 314 3787 354
rect 3721 212 3757 252
rect 3763 205 3787 245
rect 4067 226 4119 250
rect 3876 197 3913 223
rect 3876 152 3913 178
rect 3722 93 3758 133
rect 3764 86 3788 126
rect 3876 108 3913 134
rect 3876 70 3913 102
rect 3726 -15 3762 25
rect 3768 -22 3792 18
<< ntransistor >>
rect 4164 1213 4174 1215
rect 4168 1173 4178 1175
rect 4351 1152 4361 1154
rect 3621 1131 3631 1133
rect 4168 1130 4178 1132
rect 4528 1128 4538 1130
rect 4168 1122 4178 1124
rect 4355 1104 4365 1106
rect 3621 1095 3631 1097
rect 3621 1087 3631 1089
rect 4168 1086 4178 1088
rect 4532 1081 4542 1083
rect 4168 1078 4178 1080
rect 3522 1059 3532 1061
rect 4355 1061 4365 1063
rect 3621 1051 3631 1053
rect 4355 1053 4365 1055
rect 3621 1043 3631 1045
rect 4168 1042 4178 1044
rect 4532 1038 4542 1040
rect 4532 1030 4542 1032
rect 3522 1023 3532 1025
rect 3522 1015 3532 1017
rect 4355 1017 4365 1019
rect 3952 1013 3962 1015
rect 4355 1009 4365 1011
rect 3621 1000 3631 1002
rect 4532 994 4542 996
rect 4532 986 4542 988
rect 3522 979 3532 981
rect 3426 971 3436 973
rect 3522 971 3532 973
rect 4355 973 4365 975
rect 3699 941 3701 947
rect 3956 964 3966 966
rect 3426 935 3436 937
rect 3324 930 3334 932
rect 4135 963 4147 965
rect 4135 953 4147 955
rect 4532 950 4542 952
rect 3426 927 3436 929
rect 3522 928 3532 930
rect 3324 894 3334 896
rect 3426 891 3436 893
rect 4135 935 4147 937
rect 3956 921 3966 923
rect 4135 925 4147 927
rect 4304 919 4316 921
rect 3956 913 3966 915
rect 4304 909 4316 911
rect 3738 892 3740 904
rect 3748 892 3750 904
rect 3766 892 3768 904
rect 3776 892 3778 904
rect 3324 886 3334 888
rect 3699 886 3701 892
rect 4092 886 4098 888
rect 4147 886 4153 888
rect 3426 883 3436 885
rect 4304 891 4316 893
rect 3956 877 3966 879
rect 4487 889 4499 891
rect 4304 881 4316 883
rect 4487 879 4499 881
rect 3956 869 3966 871
rect 4487 861 4499 863
rect 3324 850 3334 852
rect 3324 842 3334 844
rect 3426 840 3436 842
rect 3220 833 3230 835
rect 4487 851 4499 853
rect 4261 842 4267 844
rect 4316 842 4322 844
rect 3700 809 3702 815
rect 3956 833 3966 835
rect 3123 798 3133 800
rect 3324 799 3334 801
rect 4444 812 4450 814
rect 4499 812 4505 814
rect 3220 797 3230 799
rect 3220 789 3230 791
rect 3123 762 3133 764
rect 4097 796 4117 798
rect 3944 774 3956 776
rect 3739 760 3741 772
rect 3749 760 3751 772
rect 3767 760 3769 772
rect 3777 760 3779 772
rect 3123 754 3133 756
rect 3220 753 3230 755
rect 3700 754 3702 760
rect 3944 764 3956 766
rect 4264 753 4284 755
rect 3220 745 3230 747
rect 3944 746 3956 748
rect 4446 746 4466 748
rect 3944 736 3956 738
rect 3021 725 3031 727
rect 3123 718 3133 720
rect 3123 710 3133 712
rect 3220 702 3230 704
rect 3901 697 3907 699
rect 3956 697 3962 699
rect 3021 689 3031 691
rect 3021 681 3031 683
rect 2914 668 2924 670
rect 3123 667 3133 669
rect 3703 665 3705 671
rect 3021 645 3031 647
rect 3021 637 3031 639
rect 2914 632 2924 634
rect 2914 624 2924 626
rect 3742 616 3744 628
rect 3752 616 3754 628
rect 3770 616 3772 628
rect 3780 616 3782 628
rect 3703 610 3705 616
rect 3021 594 3031 596
rect 2914 588 2924 590
rect 2914 580 2924 582
rect 4679 579 4681 599
rect 4722 581 4724 591
rect 4758 581 4760 591
rect 4766 581 4768 591
rect 4802 581 4804 591
rect 4810 581 4812 591
rect 4853 581 4855 591
rect 4891 582 4893 592
rect 3710 540 3712 546
rect 2914 537 2924 539
rect 4521 506 4621 508
rect 3749 491 3751 503
rect 3759 491 3761 503
rect 3777 491 3779 503
rect 3787 491 3789 503
rect 4333 498 4433 500
rect 3710 485 3712 491
rect 4152 488 4252 490
rect 3984 480 4084 482
rect 4523 397 4623 399
rect 4331 387 4431 389
rect 4151 377 4251 379
rect 3732 278 3734 298
rect 3743 278 3745 298
rect 3774 296 3776 306
rect 3936 269 3938 369
rect 3983 366 4083 368
rect 4016 268 4116 270
rect 4131 237 4151 239
rect 3929 208 3939 210
rect 3732 169 3734 189
rect 3743 169 3745 189
rect 3774 187 3776 197
rect 3929 165 3939 167
rect 3929 157 3939 159
rect 3929 121 3939 123
rect 3929 113 3939 115
rect 3733 50 3735 70
rect 3744 50 3746 70
rect 3775 68 3777 78
rect 3929 77 3939 79
rect 3737 -58 3739 -38
rect 3748 -58 3750 -38
rect 3779 -40 3781 -30
<< ptransistor >>
rect 4126 1213 4146 1215
rect 4121 1173 4146 1175
rect 4313 1152 4333 1154
rect 3653 1127 3678 1129
rect 4121 1128 4146 1130
rect 4490 1128 4510 1130
rect 3653 1119 3678 1121
rect 4308 1104 4333 1106
rect 3653 1089 3678 1091
rect 4121 1084 4146 1086
rect 4485 1081 4510 1083
rect 3554 1055 3579 1057
rect 4308 1059 4333 1061
rect 4121 1054 4146 1056
rect 3554 1047 3579 1049
rect 3653 1045 3678 1047
rect 4121 1046 4146 1048
rect 4485 1036 4510 1038
rect 3554 1017 3579 1019
rect 4308 1015 4333 1017
rect 3914 1013 3934 1015
rect 3653 1000 3678 1002
rect 4485 992 4510 994
rect 4308 985 4333 987
rect 4308 977 4333 979
rect 3554 973 3579 975
rect 3458 967 3483 969
rect 3699 961 3701 973
rect 3458 959 3483 961
rect 3738 945 3740 969
rect 3748 945 3750 969
rect 3909 964 3934 966
rect 3458 929 3483 931
rect 3766 939 3768 963
rect 3776 939 3778 963
rect 4076 963 4100 965
rect 4485 962 4510 964
rect 4076 953 4100 955
rect 4485 954 4510 956
rect 3356 926 3381 928
rect 3554 928 3579 930
rect 3356 918 3381 920
rect 3699 906 3701 918
rect 4070 935 4094 937
rect 4070 925 4094 927
rect 3909 919 3934 921
rect 4245 919 4269 921
rect 4245 909 4269 911
rect 3356 888 3381 890
rect 3458 885 3483 887
rect 4239 891 4263 893
rect 4066 886 4078 888
rect 4121 886 4133 888
rect 4239 881 4263 883
rect 3909 875 3934 877
rect 4428 889 4452 891
rect 4428 879 4452 881
rect 4422 861 4446 863
rect 4422 851 4446 853
rect 3356 844 3381 846
rect 3909 845 3934 847
rect 3458 840 3483 842
rect 3252 829 3277 831
rect 3700 829 3702 841
rect 4235 842 4247 844
rect 4290 842 4302 844
rect 3909 837 3934 839
rect 3252 821 3277 823
rect 3739 813 3741 837
rect 3749 813 3751 837
rect 3356 799 3381 801
rect 3767 807 3769 831
rect 3777 807 3779 831
rect 4418 812 4430 814
rect 4473 812 4485 814
rect 3155 794 3180 796
rect 3252 791 3277 793
rect 3155 786 3180 788
rect 3700 774 3702 786
rect 4039 796 4079 798
rect 3885 774 3909 776
rect 3885 764 3909 766
rect 3155 756 3180 758
rect 4206 753 4246 755
rect 3252 747 3277 749
rect 3879 746 3903 748
rect 3879 736 3903 738
rect 4388 746 4428 748
rect 3053 721 3078 723
rect 3053 713 3078 715
rect 3155 712 3180 714
rect 3252 702 3277 704
rect 3875 697 3887 699
rect 3930 697 3942 699
rect 3703 685 3705 697
rect 3053 683 3078 685
rect 3155 667 3180 669
rect 2946 664 2971 666
rect 3742 669 3744 693
rect 3752 669 3754 693
rect 2946 656 2971 658
rect 3770 663 3772 687
rect 3780 663 3782 687
rect 3053 639 3078 641
rect 3703 630 3705 642
rect 2946 626 2971 628
rect 4679 617 4681 657
rect 4726 613 4728 638
rect 4734 613 4736 638
rect 4764 613 4766 638
rect 4808 613 4810 638
rect 4853 613 4855 638
rect 3053 594 3078 596
rect 4545 591 4595 593
rect 2946 582 2971 584
rect 4891 610 4893 630
rect 3710 560 3712 572
rect 3749 544 3751 568
rect 3759 544 3761 568
rect 2946 537 2971 539
rect 3777 538 3779 562
rect 3787 538 3789 562
rect 4349 556 4399 558
rect 4175 552 4225 554
rect 3710 505 3712 517
rect 4001 529 4051 531
rect 3732 327 3734 347
rect 3743 327 3745 347
rect 3774 320 3776 340
rect 3732 218 3734 238
rect 3743 218 3745 238
rect 4073 237 4113 239
rect 3774 211 3776 231
rect 3882 208 3907 210
rect 3882 163 3907 165
rect 3882 119 3907 121
rect 3733 99 3735 119
rect 3744 99 3746 119
rect 3775 92 3777 112
rect 3882 89 3907 91
rect 3882 81 3907 83
rect 3737 -9 3739 11
rect 3748 -9 3750 11
rect 3779 -16 3781 4
<< ndiffusion >>
rect 4164 1215 4174 1216
rect 4164 1212 4174 1213
rect 4168 1175 4178 1176
rect 4168 1172 4178 1173
rect 4351 1154 4361 1155
rect 4351 1151 4361 1152
rect 3621 1133 3631 1134
rect 3621 1130 3631 1131
rect 4168 1132 4178 1133
rect 4528 1130 4538 1131
rect 4168 1129 4178 1130
rect 4168 1124 4178 1125
rect 4528 1127 4538 1128
rect 4168 1121 4178 1122
rect 4355 1106 4365 1107
rect 3621 1097 3631 1098
rect 4355 1103 4365 1104
rect 3621 1094 3631 1095
rect 3621 1089 3631 1090
rect 3621 1086 3631 1087
rect 4168 1088 4178 1089
rect 4168 1085 4178 1086
rect 4532 1083 4542 1084
rect 4168 1080 4178 1081
rect 4168 1077 4178 1078
rect 4532 1080 4542 1081
rect 3522 1061 3532 1062
rect 3522 1058 3532 1059
rect 4355 1063 4365 1064
rect 3621 1053 3631 1054
rect 4355 1060 4365 1061
rect 4355 1055 4365 1056
rect 3621 1050 3631 1051
rect 3621 1045 3631 1046
rect 3621 1042 3631 1043
rect 4355 1052 4365 1053
rect 4168 1044 4178 1045
rect 4168 1041 4178 1042
rect 4532 1040 4542 1041
rect 4532 1037 4542 1038
rect 4532 1032 4542 1033
rect 3522 1025 3532 1026
rect 4532 1029 4542 1030
rect 3522 1022 3532 1023
rect 3522 1017 3532 1018
rect 3522 1014 3532 1015
rect 4355 1019 4365 1020
rect 3952 1015 3962 1016
rect 3952 1012 3962 1013
rect 4355 1016 4365 1017
rect 4355 1011 4365 1012
rect 3621 1002 3631 1003
rect 4355 1008 4365 1009
rect 3621 999 3631 1000
rect 4532 996 4542 997
rect 4532 993 4542 994
rect 4532 988 4542 989
rect 3522 981 3532 982
rect 4532 985 4542 986
rect 3522 978 3532 979
rect 3426 973 3436 974
rect 3426 970 3436 971
rect 3522 973 3532 974
rect 3522 970 3532 971
rect 4355 975 4365 976
rect 3426 937 3436 938
rect 3698 941 3699 947
rect 3701 941 3702 947
rect 3956 966 3966 967
rect 4355 972 4365 973
rect 3324 932 3334 933
rect 3426 934 3436 935
rect 3324 929 3334 930
rect 3426 929 3436 930
rect 3522 930 3532 931
rect 3956 963 3966 964
rect 4135 965 4147 966
rect 4135 955 4147 963
rect 4135 952 4147 953
rect 4532 952 4542 953
rect 4532 949 4542 950
rect 3426 926 3436 927
rect 3522 927 3532 928
rect 3324 896 3334 897
rect 3324 893 3334 894
rect 3324 888 3334 889
rect 3426 893 3436 894
rect 4135 937 4147 938
rect 3956 923 3966 924
rect 3956 920 3966 921
rect 4135 927 4147 935
rect 4135 924 4147 925
rect 3956 915 3966 916
rect 4304 921 4316 922
rect 3956 912 3966 913
rect 4304 911 4316 919
rect 4304 908 4316 909
rect 3737 892 3738 904
rect 3740 892 3748 904
rect 3750 892 3751 904
rect 3765 892 3766 904
rect 3768 892 3776 904
rect 3778 892 3779 904
rect 4304 893 4316 894
rect 3426 890 3436 891
rect 3324 885 3334 886
rect 3426 885 3436 886
rect 3698 886 3699 892
rect 3701 886 3702 892
rect 4092 888 4098 889
rect 4147 888 4153 889
rect 3426 882 3436 883
rect 4092 885 4098 886
rect 4147 885 4153 886
rect 3956 879 3966 880
rect 3956 876 3966 877
rect 4304 883 4316 891
rect 4487 891 4499 892
rect 4487 881 4499 889
rect 4304 880 4316 881
rect 4487 878 4499 879
rect 3956 871 3966 872
rect 3956 868 3966 869
rect 4487 863 4499 864
rect 3324 852 3334 853
rect 3324 849 3334 850
rect 3324 844 3334 845
rect 3324 841 3334 842
rect 3220 835 3230 836
rect 3426 842 3436 843
rect 3426 839 3436 840
rect 3220 832 3230 833
rect 4261 844 4267 845
rect 4487 853 4499 861
rect 4487 850 4499 851
rect 4316 844 4322 845
rect 3699 809 3700 815
rect 3702 809 3703 815
rect 4261 841 4267 842
rect 4316 841 4322 842
rect 3956 835 3966 836
rect 3123 800 3133 801
rect 3123 797 3133 798
rect 3220 799 3230 800
rect 3324 801 3334 802
rect 3956 832 3966 833
rect 4444 814 4450 815
rect 4499 814 4505 815
rect 4444 811 4450 812
rect 4499 811 4505 812
rect 3324 798 3334 799
rect 3220 796 3230 797
rect 3220 791 3230 792
rect 3220 788 3230 789
rect 3123 764 3133 765
rect 3123 761 3133 762
rect 3123 756 3133 757
rect 4097 798 4117 799
rect 4097 795 4117 796
rect 3944 776 3956 777
rect 3738 760 3739 772
rect 3741 760 3749 772
rect 3751 760 3752 772
rect 3766 760 3767 772
rect 3769 760 3777 772
rect 3779 760 3780 772
rect 3944 766 3956 774
rect 3220 755 3230 756
rect 3123 753 3133 754
rect 3699 754 3700 760
rect 3702 754 3703 760
rect 3944 763 3956 764
rect 4264 755 4284 756
rect 3220 752 3230 753
rect 3220 747 3230 748
rect 3944 748 3956 749
rect 4264 752 4284 753
rect 4446 748 4466 749
rect 3220 744 3230 745
rect 3021 727 3031 728
rect 3944 738 3956 746
rect 4446 745 4466 746
rect 3944 735 3956 736
rect 3021 724 3031 725
rect 3123 720 3133 721
rect 3123 717 3133 718
rect 3123 712 3133 713
rect 3123 709 3133 710
rect 3220 704 3230 705
rect 3220 701 3230 702
rect 3901 699 3907 700
rect 3956 699 3962 700
rect 3021 691 3031 692
rect 3021 688 3031 689
rect 3021 683 3031 684
rect 3021 680 3031 681
rect 2914 670 2924 671
rect 2914 667 2924 668
rect 3123 669 3133 670
rect 3123 666 3133 667
rect 3702 665 3703 671
rect 3705 665 3706 671
rect 3901 696 3907 697
rect 3956 696 3962 697
rect 3021 647 3031 648
rect 3021 644 3031 645
rect 3021 639 3031 640
rect 2914 634 2924 635
rect 3021 636 3031 637
rect 2914 631 2924 632
rect 2914 626 2924 627
rect 2914 623 2924 624
rect 3741 616 3742 628
rect 3744 616 3752 628
rect 3754 616 3755 628
rect 3769 616 3770 628
rect 3772 616 3780 628
rect 3782 616 3783 628
rect 3702 610 3703 616
rect 3705 610 3706 616
rect 3021 596 3031 597
rect 2914 590 2924 591
rect 3021 593 3031 594
rect 2914 587 2924 588
rect 2914 582 2924 583
rect 2914 579 2924 580
rect 4678 579 4679 599
rect 4681 579 4682 599
rect 4721 581 4722 591
rect 4724 581 4725 591
rect 4757 581 4758 591
rect 4760 581 4761 591
rect 4765 581 4766 591
rect 4768 581 4769 591
rect 4801 581 4802 591
rect 4804 581 4805 591
rect 4809 581 4810 591
rect 4812 581 4813 591
rect 4852 581 4853 591
rect 4855 581 4856 591
rect 4890 582 4891 592
rect 4893 582 4894 592
rect 2914 539 2924 540
rect 3709 540 3710 546
rect 3712 540 3713 546
rect 2914 536 2924 537
rect 4521 508 4621 509
rect 4521 505 4621 506
rect 3748 491 3749 503
rect 3751 491 3759 503
rect 3761 491 3762 503
rect 3776 491 3777 503
rect 3779 491 3787 503
rect 3789 491 3790 503
rect 4333 500 4433 501
rect 4333 497 4433 498
rect 3709 485 3710 491
rect 3712 485 3713 491
rect 4152 490 4252 491
rect 4152 487 4252 488
rect 3984 482 4084 483
rect 3984 479 4084 480
rect 4523 399 4623 400
rect 4523 396 4623 397
rect 4331 389 4431 390
rect 4331 386 4431 387
rect 4151 379 4251 380
rect 4151 376 4251 377
rect 3731 278 3732 298
rect 3734 278 3743 298
rect 3745 278 3746 298
rect 3773 296 3774 306
rect 3776 296 3777 306
rect 3935 269 3936 369
rect 3938 269 3939 369
rect 3983 368 4083 369
rect 3983 365 4083 366
rect 4016 270 4116 271
rect 4016 267 4116 268
rect 4131 239 4151 240
rect 4131 236 4151 237
rect 3929 210 3939 211
rect 3929 207 3939 208
rect 3731 169 3732 189
rect 3734 169 3743 189
rect 3745 169 3746 189
rect 3773 187 3774 197
rect 3776 187 3777 197
rect 3929 167 3939 168
rect 3929 164 3939 165
rect 3929 159 3939 160
rect 3929 156 3939 157
rect 3929 123 3939 124
rect 3929 120 3939 121
rect 3929 115 3939 116
rect 3929 112 3939 113
rect 3732 50 3733 70
rect 3735 50 3744 70
rect 3746 50 3747 70
rect 3774 68 3775 78
rect 3777 68 3778 78
rect 3929 79 3939 80
rect 3929 76 3939 77
rect 3736 -58 3737 -38
rect 3739 -58 3748 -38
rect 3750 -58 3751 -38
rect 3778 -40 3779 -30
rect 3781 -40 3782 -30
<< pdiffusion >>
rect 4126 1215 4146 1216
rect 4126 1212 4146 1213
rect 4121 1175 4146 1176
rect 4121 1172 4146 1173
rect 4313 1154 4333 1155
rect 4313 1151 4333 1152
rect 4121 1130 4146 1131
rect 4490 1130 4510 1131
rect 3653 1129 3678 1130
rect 4121 1127 4146 1128
rect 3653 1126 3678 1127
rect 4490 1127 4510 1128
rect 3653 1121 3678 1122
rect 3653 1118 3678 1119
rect 4308 1106 4333 1107
rect 4308 1103 4333 1104
rect 3653 1091 3678 1092
rect 3653 1088 3678 1089
rect 4121 1086 4146 1087
rect 4121 1083 4146 1084
rect 4485 1083 4510 1084
rect 4485 1080 4510 1081
rect 4308 1061 4333 1062
rect 3554 1057 3579 1058
rect 3554 1054 3579 1055
rect 4121 1056 4146 1057
rect 4308 1058 4333 1059
rect 4121 1053 4146 1054
rect 3554 1049 3579 1050
rect 3554 1046 3579 1047
rect 4121 1048 4146 1049
rect 3653 1047 3678 1048
rect 4121 1045 4146 1046
rect 3653 1044 3678 1045
rect 4485 1038 4510 1039
rect 4485 1035 4510 1036
rect 3554 1019 3579 1020
rect 3554 1016 3579 1017
rect 3914 1015 3934 1016
rect 4308 1017 4333 1018
rect 4308 1014 4333 1015
rect 3914 1012 3934 1013
rect 3653 1002 3678 1003
rect 3653 999 3678 1000
rect 4485 994 4510 995
rect 4308 987 4333 988
rect 4485 991 4510 992
rect 4308 984 4333 985
rect 4308 979 4333 980
rect 4308 976 4333 977
rect 3554 975 3579 976
rect 3554 972 3579 973
rect 3458 969 3483 970
rect 3458 966 3483 967
rect 3458 961 3483 962
rect 3698 961 3699 973
rect 3701 961 3702 973
rect 3458 958 3483 959
rect 3737 945 3738 969
rect 3740 945 3742 969
rect 3746 945 3748 969
rect 3750 945 3751 969
rect 3909 966 3934 967
rect 4076 965 4100 966
rect 3909 963 3934 964
rect 3458 931 3483 932
rect 3765 939 3766 963
rect 3768 939 3770 963
rect 3774 939 3776 963
rect 3778 939 3779 963
rect 4076 961 4100 963
rect 4485 964 4510 965
rect 4076 955 4100 957
rect 4485 961 4510 962
rect 4485 956 4510 957
rect 4076 952 4100 953
rect 4485 953 4510 954
rect 3554 930 3579 931
rect 3356 928 3381 929
rect 3458 928 3483 929
rect 3356 925 3381 926
rect 3554 927 3579 928
rect 3356 920 3381 921
rect 3356 917 3381 918
rect 3698 906 3699 918
rect 3701 906 3702 918
rect 4070 937 4094 938
rect 4070 933 4094 935
rect 4070 927 4094 929
rect 4070 924 4094 925
rect 3909 921 3934 922
rect 3909 918 3934 919
rect 4245 921 4269 922
rect 4245 917 4269 919
rect 4245 911 4269 913
rect 4245 908 4269 909
rect 4239 893 4263 894
rect 3356 890 3381 891
rect 3356 887 3381 888
rect 3458 887 3483 888
rect 4066 888 4078 889
rect 4121 888 4133 889
rect 4239 889 4263 891
rect 3458 884 3483 885
rect 4066 885 4078 886
rect 4121 885 4133 886
rect 4428 891 4452 892
rect 4239 883 4263 885
rect 4239 880 4263 881
rect 3909 877 3934 878
rect 3909 874 3934 875
rect 4428 887 4452 889
rect 4428 881 4452 883
rect 4428 878 4452 879
rect 4422 863 4446 864
rect 4422 859 4446 861
rect 4422 853 4446 855
rect 4422 850 4446 851
rect 3909 847 3934 848
rect 3356 846 3381 847
rect 3356 843 3381 844
rect 3909 844 3934 845
rect 3458 842 3483 843
rect 3458 839 3483 840
rect 3252 831 3277 832
rect 3699 829 3700 841
rect 3702 829 3703 841
rect 4235 844 4247 845
rect 4290 844 4302 845
rect 4235 841 4247 842
rect 3909 839 3934 840
rect 3252 828 3277 829
rect 3252 823 3277 824
rect 3252 820 3277 821
rect 3738 813 3739 837
rect 3741 813 3743 837
rect 3747 813 3749 837
rect 3751 813 3752 837
rect 3909 836 3934 837
rect 4290 841 4302 842
rect 3356 801 3381 802
rect 3766 807 3767 831
rect 3769 807 3771 831
rect 3775 807 3777 831
rect 3779 807 3780 831
rect 4418 814 4430 815
rect 4473 814 4485 815
rect 4418 811 4430 812
rect 4473 811 4485 812
rect 3155 796 3180 797
rect 3155 793 3180 794
rect 3356 798 3381 799
rect 3252 793 3277 794
rect 3252 790 3277 791
rect 3155 788 3180 789
rect 3155 785 3180 786
rect 3699 774 3700 786
rect 3702 774 3703 786
rect 4039 798 4079 799
rect 4039 795 4079 796
rect 3885 776 3909 777
rect 3885 772 3909 774
rect 3885 766 3909 768
rect 3885 763 3909 764
rect 3155 758 3180 759
rect 3155 755 3180 756
rect 4206 755 4246 756
rect 3252 749 3277 750
rect 3879 748 3903 749
rect 4206 752 4246 753
rect 4388 748 4428 749
rect 3252 746 3277 747
rect 3879 744 3903 746
rect 3879 738 3903 740
rect 3879 735 3903 736
rect 4388 745 4428 746
rect 3053 723 3078 724
rect 3053 720 3078 721
rect 3053 715 3078 716
rect 3053 712 3078 713
rect 3155 714 3180 715
rect 3155 711 3180 712
rect 3252 704 3277 705
rect 3252 701 3277 702
rect 3875 699 3887 700
rect 3930 699 3942 700
rect 3053 685 3078 686
rect 3702 685 3703 697
rect 3705 685 3706 697
rect 3875 696 3887 697
rect 3053 682 3078 683
rect 3155 669 3180 670
rect 2946 666 2971 667
rect 2946 663 2971 664
rect 3155 666 3180 667
rect 3741 669 3742 693
rect 3744 669 3746 693
rect 3750 669 3752 693
rect 3754 669 3755 693
rect 3930 696 3942 697
rect 2946 658 2971 659
rect 2946 655 2971 656
rect 3769 663 3770 687
rect 3772 663 3774 687
rect 3778 663 3780 687
rect 3782 663 3783 687
rect 3053 641 3078 642
rect 3053 638 3078 639
rect 3702 630 3703 642
rect 3705 630 3706 642
rect 2946 628 2971 629
rect 2946 625 2971 626
rect 4678 617 4679 657
rect 4681 617 4682 657
rect 4725 613 4726 638
rect 4728 613 4729 638
rect 4733 613 4734 638
rect 4736 613 4737 638
rect 4763 613 4764 638
rect 4766 613 4767 638
rect 4807 613 4808 638
rect 4810 613 4811 638
rect 4852 613 4853 638
rect 4855 613 4856 638
rect 3053 596 3078 597
rect 3053 593 3078 594
rect 4545 593 4595 594
rect 4545 590 4595 591
rect 2946 584 2971 585
rect 2946 581 2971 582
rect 4890 610 4891 630
rect 4893 610 4894 630
rect 3709 560 3710 572
rect 3712 560 3713 572
rect 3748 544 3749 568
rect 3751 544 3753 568
rect 3757 544 3759 568
rect 3761 544 3762 568
rect 2946 539 2971 540
rect 2946 536 2971 537
rect 3776 538 3777 562
rect 3779 538 3781 562
rect 3785 538 3787 562
rect 3789 538 3790 562
rect 4175 554 4225 555
rect 4349 558 4399 559
rect 4349 555 4399 556
rect 4175 551 4225 552
rect 3709 505 3710 517
rect 3712 505 3713 517
rect 4001 531 4051 532
rect 4001 528 4051 529
rect 3731 327 3732 347
rect 3734 327 3738 347
rect 3742 327 3743 347
rect 3745 327 3746 347
rect 3773 320 3774 340
rect 3776 320 3777 340
rect 4073 239 4113 240
rect 3731 218 3732 238
rect 3734 218 3738 238
rect 3742 218 3743 238
rect 3745 218 3746 238
rect 4073 236 4113 237
rect 3773 211 3774 231
rect 3776 211 3777 231
rect 3882 210 3907 211
rect 3882 207 3907 208
rect 3882 165 3907 166
rect 3882 162 3907 163
rect 3882 121 3907 122
rect 3732 99 3733 119
rect 3735 99 3739 119
rect 3743 99 3744 119
rect 3746 99 3747 119
rect 3882 118 3907 119
rect 3774 92 3775 112
rect 3777 92 3778 112
rect 3882 91 3907 92
rect 3882 88 3907 89
rect 3882 83 3907 84
rect 3882 80 3907 81
rect 3736 -9 3737 11
rect 3739 -9 3743 11
rect 3747 -9 3748 11
rect 3750 -9 3751 11
rect 3778 -16 3779 4
rect 3781 -16 3782 4
<< ndcontact >>
rect 4164 1216 4174 1220
rect 4164 1208 4174 1212
rect 4168 1176 4178 1180
rect 4168 1168 4178 1172
rect 4351 1155 4361 1159
rect 4351 1147 4361 1151
rect 3621 1134 3631 1138
rect 3621 1126 3631 1130
rect 4168 1133 4178 1137
rect 4528 1131 4538 1135
rect 4168 1125 4178 1129
rect 4528 1123 4538 1127
rect 4168 1117 4178 1121
rect 4355 1107 4365 1111
rect 3621 1098 3631 1102
rect 4355 1099 4365 1103
rect 3621 1090 3631 1094
rect 3621 1082 3631 1086
rect 4168 1089 4178 1093
rect 4168 1081 4178 1085
rect 4532 1084 4542 1088
rect 4168 1073 4178 1077
rect 4532 1076 4542 1080
rect 3522 1062 3532 1066
rect 3522 1054 3532 1058
rect 4355 1064 4365 1068
rect 3621 1054 3631 1058
rect 4355 1056 4365 1060
rect 3621 1046 3631 1050
rect 3621 1038 3631 1042
rect 4168 1045 4178 1049
rect 4355 1048 4365 1052
rect 4168 1037 4178 1041
rect 4532 1041 4542 1045
rect 4532 1033 4542 1037
rect 3522 1026 3532 1030
rect 4532 1025 4542 1029
rect 3522 1018 3532 1022
rect 3522 1010 3532 1014
rect 3952 1016 3962 1020
rect 4355 1020 4365 1024
rect 3952 1008 3962 1012
rect 4355 1012 4365 1016
rect 3621 1003 3631 1007
rect 4355 1004 4365 1008
rect 3621 995 3631 999
rect 4532 997 4542 1001
rect 4532 989 4542 993
rect 3522 982 3532 986
rect 4532 981 4542 985
rect 3426 974 3436 978
rect 3522 974 3532 978
rect 3426 966 3436 970
rect 3522 966 3532 970
rect 4355 976 4365 980
rect 3426 938 3436 942
rect 3694 941 3698 947
rect 3702 941 3706 947
rect 3956 967 3966 971
rect 4135 966 4147 970
rect 4355 968 4365 972
rect 3324 933 3334 937
rect 3324 925 3334 929
rect 3426 930 3436 934
rect 3522 931 3532 935
rect 3956 959 3966 963
rect 4135 948 4147 952
rect 4532 953 4542 957
rect 4532 945 4542 949
rect 3426 922 3436 926
rect 3522 923 3532 927
rect 3324 897 3334 901
rect 3324 889 3334 893
rect 3426 894 3436 898
rect 4135 938 4147 942
rect 3956 924 3966 928
rect 4135 920 4147 924
rect 4304 922 4316 926
rect 3956 916 3966 920
rect 3956 908 3966 912
rect 4304 904 4316 908
rect 3733 892 3737 904
rect 3751 892 3755 904
rect 3761 892 3765 904
rect 3779 892 3783 904
rect 4304 894 4316 898
rect 3324 881 3334 885
rect 3426 886 3436 890
rect 3694 886 3698 892
rect 3702 886 3706 892
rect 4092 889 4098 893
rect 4147 889 4153 893
rect 3426 878 3436 882
rect 3956 880 3966 884
rect 4092 881 4098 885
rect 4147 881 4153 885
rect 4487 892 4499 896
rect 4304 876 4316 880
rect 3956 872 3966 876
rect 4487 874 4499 878
rect 3956 864 3966 868
rect 4487 864 4499 868
rect 3324 853 3334 857
rect 3324 845 3334 849
rect 3220 836 3230 840
rect 3324 837 3334 841
rect 3426 843 3436 847
rect 3220 828 3230 832
rect 3426 835 3436 839
rect 4261 845 4267 849
rect 4316 845 4322 849
rect 4487 846 4499 850
rect 3695 809 3699 815
rect 3703 809 3707 815
rect 3956 836 3966 840
rect 4261 837 4267 841
rect 4316 837 4322 841
rect 3123 801 3133 805
rect 3123 793 3133 797
rect 3220 800 3230 804
rect 3324 802 3334 806
rect 3956 828 3966 832
rect 4444 815 4450 819
rect 4499 815 4505 819
rect 4444 807 4450 811
rect 4499 807 4505 811
rect 3220 792 3230 796
rect 3324 794 3334 798
rect 3220 784 3230 788
rect 3123 765 3133 769
rect 3123 757 3133 761
rect 4097 799 4117 803
rect 4097 791 4117 795
rect 3944 777 3956 781
rect 3734 760 3738 772
rect 3752 760 3756 772
rect 3762 760 3766 772
rect 3780 760 3784 772
rect 3220 756 3230 760
rect 3123 749 3133 753
rect 3695 754 3699 760
rect 3703 754 3707 760
rect 3944 759 3956 763
rect 4264 756 4284 760
rect 3220 748 3230 752
rect 3944 749 3956 753
rect 4264 748 4284 752
rect 4446 749 4466 753
rect 3220 740 3230 744
rect 3021 728 3031 732
rect 4446 741 4466 745
rect 3944 731 3956 735
rect 3021 720 3031 724
rect 3123 721 3133 725
rect 3123 713 3133 717
rect 3123 705 3133 709
rect 3220 705 3230 709
rect 3220 697 3230 701
rect 3901 700 3907 704
rect 3956 700 3962 704
rect 3021 692 3031 696
rect 3021 684 3031 688
rect 3021 676 3031 680
rect 2914 671 2924 675
rect 2914 663 2924 667
rect 3123 670 3133 674
rect 3123 662 3133 666
rect 3698 665 3702 671
rect 3706 665 3710 671
rect 3901 692 3907 696
rect 3956 692 3962 696
rect 3021 648 3031 652
rect 3021 640 3031 644
rect 2914 635 2924 639
rect 2914 627 2924 631
rect 3021 632 3031 636
rect 2914 619 2924 623
rect 3737 616 3741 628
rect 3755 616 3759 628
rect 3765 616 3769 628
rect 3783 616 3787 628
rect 3698 610 3702 616
rect 3706 610 3710 616
rect 3021 597 3031 601
rect 2914 591 2924 595
rect 3021 589 3031 593
rect 2914 583 2924 587
rect 2914 575 2924 579
rect 4674 579 4678 599
rect 4682 579 4686 599
rect 4717 581 4721 591
rect 4725 581 4729 591
rect 4753 581 4757 591
rect 4761 581 4765 591
rect 4769 581 4773 591
rect 4797 581 4801 591
rect 4805 581 4809 591
rect 4813 581 4817 591
rect 4848 581 4852 591
rect 4856 581 4860 591
rect 4886 582 4890 592
rect 4894 582 4898 592
rect 2914 540 2924 544
rect 3705 540 3709 546
rect 3713 540 3717 546
rect 2914 532 2924 536
rect 4521 509 4621 513
rect 3744 491 3748 503
rect 3762 491 3766 503
rect 3772 491 3776 503
rect 3790 491 3794 503
rect 4333 501 4433 505
rect 4521 501 4621 505
rect 3705 485 3709 491
rect 3713 485 3717 491
rect 4152 491 4252 495
rect 4333 493 4433 497
rect 3984 483 4084 487
rect 4152 483 4252 487
rect 3984 475 4084 479
rect 4523 400 4623 404
rect 4331 390 4431 394
rect 4523 392 4623 396
rect 4151 380 4251 384
rect 4331 382 4431 386
rect 3727 278 3731 298
rect 3746 278 3750 298
rect 3769 296 3773 306
rect 3777 296 3781 306
rect 3931 269 3935 369
rect 3939 269 3943 369
rect 3983 369 4083 373
rect 4151 372 4251 376
rect 3983 361 4083 365
rect 4016 271 4116 275
rect 4016 263 4116 267
rect 4131 240 4151 244
rect 4131 232 4151 236
rect 3929 211 3939 215
rect 3929 203 3939 207
rect 3727 169 3731 189
rect 3746 169 3750 189
rect 3769 187 3773 197
rect 3777 187 3781 197
rect 3929 168 3939 172
rect 3929 160 3939 164
rect 3929 152 3939 156
rect 3929 124 3939 128
rect 3929 116 3939 120
rect 3929 108 3939 112
rect 3728 50 3732 70
rect 3747 50 3751 70
rect 3770 68 3774 78
rect 3778 68 3782 78
rect 3929 80 3939 84
rect 3929 72 3939 76
rect 3732 -58 3736 -38
rect 3751 -58 3755 -38
rect 3774 -40 3778 -30
rect 3782 -40 3786 -30
<< pdcontact >>
rect 4126 1216 4146 1220
rect 4126 1208 4146 1212
rect 4121 1176 4146 1180
rect 4121 1168 4146 1172
rect 4313 1155 4333 1159
rect 4313 1147 4333 1151
rect 3653 1130 3678 1134
rect 4121 1131 4146 1135
rect 4490 1131 4510 1135
rect 3653 1122 3678 1126
rect 4121 1123 4146 1127
rect 4490 1123 4510 1127
rect 3653 1114 3678 1118
rect 4308 1107 4333 1111
rect 4308 1099 4333 1103
rect 3653 1092 3678 1096
rect 3653 1084 3678 1088
rect 4121 1087 4146 1091
rect 4121 1079 4146 1083
rect 4485 1084 4510 1088
rect 4485 1076 4510 1080
rect 3554 1058 3579 1062
rect 4308 1062 4333 1066
rect 3554 1050 3579 1054
rect 4121 1057 4146 1061
rect 4308 1054 4333 1058
rect 3554 1042 3579 1046
rect 3653 1048 3678 1052
rect 4121 1049 4146 1053
rect 3653 1040 3678 1044
rect 4121 1041 4146 1045
rect 4485 1039 4510 1043
rect 4485 1031 4510 1035
rect 3554 1020 3579 1024
rect 3554 1012 3579 1016
rect 3914 1016 3934 1020
rect 4308 1018 4333 1022
rect 3914 1008 3934 1012
rect 4308 1010 4333 1014
rect 3653 1003 3678 1007
rect 3653 995 3678 999
rect 4485 995 4510 999
rect 4308 988 4333 992
rect 4485 987 4510 991
rect 4308 980 4333 984
rect 3458 970 3483 974
rect 3554 976 3579 980
rect 3554 968 3579 972
rect 3458 962 3483 966
rect 3694 961 3698 973
rect 3702 961 3706 973
rect 4308 972 4333 976
rect 3458 954 3483 958
rect 3733 945 3737 969
rect 3742 945 3746 969
rect 3751 945 3755 969
rect 3909 967 3934 971
rect 4076 966 4100 970
rect 3356 929 3381 933
rect 3458 932 3483 936
rect 3554 931 3579 935
rect 3761 939 3765 963
rect 3770 939 3774 963
rect 3779 939 3783 963
rect 3909 959 3934 963
rect 4485 965 4510 969
rect 4076 957 4100 961
rect 4485 957 4510 961
rect 4076 948 4100 952
rect 4485 949 4510 953
rect 3356 921 3381 925
rect 3458 924 3483 928
rect 3554 923 3579 927
rect 3356 913 3381 917
rect 3694 906 3698 918
rect 3702 906 3706 918
rect 3356 891 3381 895
rect 4070 938 4094 942
rect 4070 929 4094 933
rect 3909 922 3934 926
rect 3909 914 3934 918
rect 4070 920 4094 924
rect 4245 922 4269 926
rect 4245 913 4269 917
rect 4245 904 4269 908
rect 4239 894 4263 898
rect 3356 883 3381 887
rect 3458 888 3483 892
rect 4066 889 4078 893
rect 4121 889 4133 893
rect 3458 880 3483 884
rect 3909 878 3934 882
rect 4066 881 4078 885
rect 4121 881 4133 885
rect 4239 885 4263 889
rect 4428 892 4452 896
rect 3909 870 3934 874
rect 4239 876 4263 880
rect 4428 883 4452 887
rect 4428 874 4452 878
rect 4422 864 4446 868
rect 4422 855 4446 859
rect 3356 847 3381 851
rect 3909 848 3934 852
rect 3356 839 3381 843
rect 3458 843 3483 847
rect 3252 832 3277 836
rect 3458 835 3483 839
rect 3695 829 3699 841
rect 3703 829 3707 841
rect 3909 840 3934 844
rect 4235 845 4247 849
rect 4290 845 4302 849
rect 4422 846 4446 850
rect 3252 824 3277 828
rect 3252 816 3277 820
rect 3734 813 3738 837
rect 3743 813 3747 837
rect 3752 813 3756 837
rect 3909 832 3934 836
rect 4235 837 4247 841
rect 4290 837 4302 841
rect 3155 797 3180 801
rect 3356 802 3381 806
rect 3762 807 3766 831
rect 3771 807 3775 831
rect 3780 807 3784 831
rect 4418 815 4430 819
rect 4473 815 4485 819
rect 4418 807 4430 811
rect 4473 807 4485 811
rect 3155 789 3180 793
rect 3252 794 3277 798
rect 3356 794 3381 798
rect 3155 781 3180 785
rect 3252 786 3277 790
rect 3695 774 3699 786
rect 3703 774 3707 786
rect 3155 759 3180 763
rect 4039 799 4079 803
rect 4039 791 4079 795
rect 3885 777 3909 781
rect 3885 768 3909 772
rect 3155 751 3180 755
rect 3885 759 3909 763
rect 4206 756 4246 760
rect 3252 750 3277 754
rect 3879 749 3903 753
rect 4206 748 4246 752
rect 4388 749 4428 753
rect 3252 742 3277 746
rect 3879 740 3903 744
rect 3879 731 3903 735
rect 4388 741 4428 745
rect 3053 724 3078 728
rect 3053 716 3078 720
rect 3155 715 3180 719
rect 3053 708 3078 712
rect 3155 707 3180 711
rect 3252 705 3277 709
rect 3252 697 3277 701
rect 3875 700 3887 704
rect 3930 700 3942 704
rect 3053 686 3078 690
rect 3698 685 3702 697
rect 3706 685 3710 697
rect 3053 678 3078 682
rect 2946 667 2971 671
rect 3155 670 3180 674
rect 2946 659 2971 663
rect 3155 662 3180 666
rect 3737 669 3741 693
rect 3746 669 3750 693
rect 3755 669 3759 693
rect 3875 692 3887 696
rect 3930 692 3942 696
rect 3765 663 3769 687
rect 3774 663 3778 687
rect 3783 663 3787 687
rect 2946 651 2971 655
rect 3053 642 3078 646
rect 2946 629 2971 633
rect 3053 634 3078 638
rect 3698 630 3702 642
rect 3706 630 3710 642
rect 2946 621 2971 625
rect 4674 617 4678 657
rect 4682 617 4686 657
rect 3053 597 3078 601
rect 4721 613 4725 638
rect 4729 613 4733 638
rect 4737 613 4741 638
rect 4759 613 4763 638
rect 4767 613 4771 638
rect 4803 613 4807 638
rect 4811 613 4815 638
rect 4848 613 4852 638
rect 4856 613 4860 638
rect 4545 594 4595 598
rect 3053 589 3078 593
rect 2946 585 2971 589
rect 4545 586 4595 590
rect 2946 577 2971 581
rect 4886 610 4890 630
rect 4894 610 4898 630
rect 3705 560 3709 572
rect 3713 560 3717 572
rect 2946 540 2971 544
rect 3744 544 3748 568
rect 3753 544 3757 568
rect 3762 544 3766 568
rect 2946 532 2971 536
rect 3772 538 3776 562
rect 3781 538 3785 562
rect 3790 538 3794 562
rect 4175 555 4225 559
rect 4349 559 4399 563
rect 4349 551 4399 555
rect 4175 547 4225 551
rect 3705 505 3709 517
rect 3713 505 3717 517
rect 4001 532 4051 536
rect 4001 524 4051 528
rect 3727 327 3731 347
rect 3738 327 3742 347
rect 3746 327 3750 347
rect 3769 320 3773 340
rect 3777 320 3781 340
rect 4073 240 4113 244
rect 3727 218 3731 238
rect 3738 218 3742 238
rect 3746 218 3750 238
rect 4073 232 4113 236
rect 3769 211 3773 231
rect 3777 211 3781 231
rect 3882 211 3907 215
rect 3882 203 3907 207
rect 3882 166 3907 170
rect 3882 158 3907 162
rect 3882 122 3907 126
rect 3728 99 3732 119
rect 3739 99 3743 119
rect 3747 99 3751 119
rect 3882 114 3907 118
rect 3770 92 3774 112
rect 3778 92 3782 112
rect 3882 92 3907 96
rect 3882 84 3907 88
rect 3882 76 3907 80
rect 3732 -9 3736 11
rect 3743 -9 3747 11
rect 3751 -9 3755 11
rect 3774 -16 3778 4
rect 3782 -16 3786 4
<< psubstratepcontact >>
rect 3783 287 3788 291
rect 3783 178 3788 182
rect 3784 59 3789 63
rect 3788 -49 3793 -45
<< nsubstratencontact >>
rect 4116 1203 4120 1207
rect 4303 1142 4307 1146
rect 4480 1118 4484 1122
rect 3904 1003 3908 1007
rect 4029 786 4033 790
rect 4196 743 4200 747
rect 4378 736 4382 740
rect 4669 663 4673 667
rect 4534 599 4539 603
rect 4881 636 4885 640
rect 4338 564 4343 568
rect 4164 560 4169 564
rect 3990 537 3995 541
rect 3727 352 3731 358
rect 3779 347 3783 351
rect 3727 243 3731 249
rect 3779 238 3783 242
rect 4063 227 4067 231
rect 3728 124 3732 130
rect 3780 119 3784 123
rect 3732 16 3736 22
rect 3784 11 3788 15
<< polysilicon >>
rect 4123 1213 4126 1215
rect 4146 1213 4164 1215
rect 4174 1213 4178 1215
rect 4118 1173 4121 1175
rect 4146 1173 4168 1175
rect 4178 1173 4181 1175
rect 4310 1152 4313 1154
rect 4333 1152 4351 1154
rect 4361 1152 4365 1154
rect 3642 1133 3646 1134
rect 3618 1131 3621 1133
rect 3631 1131 3646 1133
rect 3642 1129 3646 1131
rect 4159 1130 4168 1132
rect 4178 1130 4181 1132
rect 3642 1127 3653 1129
rect 3678 1127 3681 1129
rect 4118 1128 4121 1130
rect 4146 1128 4156 1130
rect 4154 1124 4156 1128
rect 4487 1128 4490 1130
rect 4510 1128 4528 1130
rect 4538 1128 4542 1130
rect 4154 1122 4168 1124
rect 4178 1122 4181 1124
rect 3634 1119 3653 1121
rect 3678 1119 3681 1121
rect 4305 1104 4308 1106
rect 4333 1104 4355 1106
rect 4365 1104 4368 1106
rect 3618 1095 3621 1097
rect 3631 1095 3645 1097
rect 3643 1091 3645 1095
rect 3643 1089 3653 1091
rect 3678 1089 3681 1091
rect 3618 1087 3621 1089
rect 3631 1087 3640 1089
rect 4159 1086 4168 1088
rect 4178 1086 4181 1088
rect 4118 1084 4121 1086
rect 4146 1084 4156 1086
rect 4154 1080 4156 1084
rect 4482 1081 4485 1083
rect 4510 1081 4532 1083
rect 4542 1081 4545 1083
rect 4154 1078 4168 1080
rect 4178 1078 4181 1080
rect 3543 1061 3547 1062
rect 3519 1059 3522 1061
rect 3532 1059 3547 1061
rect 3543 1057 3547 1059
rect 4346 1061 4355 1063
rect 4365 1061 4368 1063
rect 3543 1055 3554 1057
rect 3579 1055 3582 1057
rect 4305 1059 4308 1061
rect 4333 1059 4343 1061
rect 4118 1054 4121 1056
rect 4146 1054 4165 1056
rect 4341 1055 4343 1059
rect 3618 1051 3621 1053
rect 3631 1051 3645 1053
rect 3535 1047 3554 1049
rect 3579 1047 3582 1049
rect 3643 1047 3645 1051
rect 4341 1053 4355 1055
rect 4365 1053 4368 1055
rect 3643 1045 3653 1047
rect 3678 1045 3681 1047
rect 4118 1046 4121 1048
rect 4146 1046 4157 1048
rect 3618 1043 3621 1045
rect 3631 1043 3640 1045
rect 4153 1044 4157 1046
rect 4153 1042 4168 1044
rect 4178 1042 4181 1044
rect 4153 1041 4157 1042
rect 4523 1038 4532 1040
rect 4542 1038 4545 1040
rect 4482 1036 4485 1038
rect 4510 1036 4520 1038
rect 4518 1032 4520 1036
rect 4518 1030 4532 1032
rect 4542 1030 4545 1032
rect 3519 1023 3522 1025
rect 3532 1023 3546 1025
rect 3544 1019 3546 1023
rect 3544 1017 3554 1019
rect 3579 1017 3582 1019
rect 3519 1015 3522 1017
rect 3532 1015 3541 1017
rect 4346 1017 4355 1019
rect 4365 1017 4368 1019
rect 4305 1015 4308 1017
rect 4333 1015 4343 1017
rect 3911 1013 3914 1015
rect 3934 1013 3952 1015
rect 3962 1013 3966 1015
rect 4341 1011 4343 1015
rect 4341 1009 4355 1011
rect 4365 1009 4368 1011
rect 3618 1000 3621 1002
rect 3631 1000 3653 1002
rect 3678 1000 3681 1002
rect 4523 994 4532 996
rect 4542 994 4545 996
rect 4482 992 4485 994
rect 4510 992 4520 994
rect 4518 988 4520 992
rect 4305 985 4308 987
rect 4333 985 4352 987
rect 4518 986 4532 988
rect 4542 986 4545 988
rect 3519 979 3522 981
rect 3532 979 3546 981
rect 3447 973 3451 974
rect 3423 971 3426 973
rect 3436 971 3451 973
rect 3447 969 3451 971
rect 3544 975 3546 979
rect 4305 977 4308 979
rect 4333 977 4344 979
rect 3544 973 3554 975
rect 3579 973 3582 975
rect 3699 973 3701 976
rect 3519 971 3522 973
rect 3532 971 3541 973
rect 3447 967 3458 969
rect 3483 967 3486 969
rect 4340 975 4344 977
rect 4340 973 4355 975
rect 4365 973 4368 975
rect 4340 972 4344 973
rect 3738 969 3740 972
rect 3748 969 3750 972
rect 3439 959 3458 961
rect 3483 959 3486 961
rect 3699 947 3701 961
rect 3766 963 3768 966
rect 3776 963 3778 966
rect 3906 964 3909 966
rect 3934 964 3956 966
rect 3966 964 3969 966
rect 3699 938 3701 941
rect 3423 935 3426 937
rect 3436 935 3450 937
rect 3738 936 3740 945
rect 3345 932 3349 933
rect 3321 930 3324 932
rect 3334 930 3349 932
rect 3345 928 3349 930
rect 3448 931 3450 935
rect 3448 929 3458 931
rect 3483 929 3486 931
rect 3748 935 3750 945
rect 4073 963 4076 965
rect 4100 963 4122 965
rect 4126 963 4135 965
rect 4147 963 4150 965
rect 4482 962 4485 964
rect 4510 962 4529 964
rect 4073 953 4076 955
rect 4100 953 4111 955
rect 4115 953 4135 955
rect 4147 953 4150 955
rect 4482 954 4485 956
rect 4510 954 4521 956
rect 4517 952 4521 954
rect 4517 950 4532 952
rect 4542 950 4545 952
rect 4517 949 4521 950
rect 3345 926 3356 928
rect 3381 926 3384 928
rect 3423 927 3426 929
rect 3436 927 3445 929
rect 3519 928 3522 930
rect 3532 928 3554 930
rect 3579 928 3582 930
rect 3337 918 3356 920
rect 3381 918 3384 920
rect 3699 918 3701 921
rect 3321 894 3324 896
rect 3334 894 3348 896
rect 3346 890 3348 894
rect 3423 891 3426 893
rect 3436 891 3450 893
rect 3699 892 3701 906
rect 3738 904 3740 931
rect 3748 904 3750 930
rect 3766 928 3768 939
rect 3766 904 3768 924
rect 3776 917 3778 939
rect 4067 935 4070 937
rect 4094 935 4104 937
rect 4109 935 4135 937
rect 4147 935 4150 937
rect 4067 925 4070 927
rect 4094 925 4103 927
rect 3947 921 3956 923
rect 3966 921 3969 923
rect 3906 919 3909 921
rect 3934 919 3944 921
rect 3942 915 3944 919
rect 4108 925 4135 927
rect 4147 925 4150 927
rect 4242 919 4245 921
rect 4269 919 4291 921
rect 4295 919 4304 921
rect 4316 919 4319 921
rect 3942 913 3956 915
rect 3966 913 3969 915
rect 3776 904 3778 913
rect 4242 909 4245 911
rect 4269 909 4280 911
rect 4284 909 4304 911
rect 4316 909 4319 911
rect 3346 888 3356 890
rect 3381 888 3384 890
rect 3321 886 3324 888
rect 3334 886 3343 888
rect 3448 887 3450 891
rect 3448 885 3458 887
rect 3483 885 3486 887
rect 3738 889 3740 892
rect 3748 889 3750 892
rect 3766 889 3768 892
rect 3776 889 3778 892
rect 4236 891 4239 893
rect 4263 891 4273 893
rect 4063 886 4066 888
rect 4078 886 4092 888
rect 4098 886 4101 888
rect 4118 886 4121 888
rect 4133 886 4147 888
rect 4153 886 4156 888
rect 3423 883 3426 885
rect 3436 883 3445 885
rect 3699 883 3701 886
rect 4278 891 4304 893
rect 4316 891 4319 893
rect 4236 881 4239 883
rect 4263 881 4272 883
rect 3947 877 3956 879
rect 3966 877 3969 879
rect 3906 875 3909 877
rect 3934 875 3944 877
rect 3942 871 3944 875
rect 4425 889 4428 891
rect 4452 889 4474 891
rect 4478 889 4487 891
rect 4499 889 4502 891
rect 4277 881 4304 883
rect 4316 881 4319 883
rect 4425 879 4428 881
rect 4452 879 4463 881
rect 4467 879 4487 881
rect 4499 879 4502 881
rect 3942 869 3956 871
rect 3966 869 3969 871
rect 4419 861 4422 863
rect 4446 861 4456 863
rect 4461 861 4487 863
rect 4499 861 4502 863
rect 3321 850 3324 852
rect 3334 850 3348 852
rect 3346 846 3348 850
rect 4419 851 4422 853
rect 4446 851 4455 853
rect 3346 844 3356 846
rect 3381 844 3384 846
rect 3321 842 3324 844
rect 3334 842 3343 844
rect 3906 845 3909 847
rect 3934 845 3953 847
rect 3423 840 3426 842
rect 3436 840 3458 842
rect 3483 840 3486 842
rect 3700 841 3702 844
rect 3241 835 3245 836
rect 3217 833 3220 835
rect 3230 833 3245 835
rect 3241 831 3245 833
rect 3241 829 3252 831
rect 3277 829 3280 831
rect 4460 851 4487 853
rect 4499 851 4502 853
rect 4232 842 4235 844
rect 4247 842 4261 844
rect 4267 842 4270 844
rect 4287 842 4290 844
rect 4302 842 4316 844
rect 4322 842 4325 844
rect 3739 837 3741 840
rect 3749 837 3751 840
rect 3906 837 3909 839
rect 3934 837 3945 839
rect 3233 821 3252 823
rect 3277 821 3280 823
rect 3700 815 3702 829
rect 3767 831 3769 834
rect 3777 831 3779 834
rect 3941 835 3945 837
rect 3941 833 3956 835
rect 3966 833 3969 835
rect 3941 832 3945 833
rect 3700 806 3702 809
rect 3144 800 3148 801
rect 3120 798 3123 800
rect 3133 798 3148 800
rect 3144 796 3148 798
rect 3739 804 3741 813
rect 3321 799 3324 801
rect 3334 799 3356 801
rect 3381 799 3384 801
rect 3749 803 3751 813
rect 4415 812 4418 814
rect 4430 812 4444 814
rect 4450 812 4453 814
rect 4470 812 4473 814
rect 4485 812 4499 814
rect 4505 812 4508 814
rect 3217 797 3220 799
rect 3230 797 3244 799
rect 3144 794 3155 796
rect 3180 794 3183 796
rect 3242 793 3244 797
rect 3242 791 3252 793
rect 3277 791 3280 793
rect 3217 789 3220 791
rect 3230 789 3239 791
rect 3136 786 3155 788
rect 3180 786 3183 788
rect 3700 786 3702 789
rect 3120 762 3123 764
rect 3133 762 3147 764
rect 3145 758 3147 762
rect 3700 760 3702 774
rect 3739 772 3741 799
rect 3749 772 3751 798
rect 3767 796 3769 807
rect 3767 772 3769 792
rect 3777 785 3779 807
rect 4036 796 4039 798
rect 4079 796 4097 798
rect 4117 796 4121 798
rect 3777 772 3779 781
rect 3882 774 3885 776
rect 3909 774 3931 776
rect 3935 774 3944 776
rect 3956 774 3959 776
rect 3882 764 3885 766
rect 3909 764 3920 766
rect 3145 756 3155 758
rect 3180 756 3183 758
rect 3120 754 3123 756
rect 3133 754 3142 756
rect 3217 753 3220 755
rect 3230 753 3244 755
rect 3739 757 3741 760
rect 3749 757 3751 760
rect 3767 757 3769 760
rect 3777 757 3779 760
rect 3924 764 3944 766
rect 3956 764 3959 766
rect 3242 749 3244 753
rect 3700 751 3702 754
rect 4203 753 4206 755
rect 4246 753 4264 755
rect 4284 753 4288 755
rect 3242 747 3252 749
rect 3277 747 3280 749
rect 3217 745 3220 747
rect 3230 745 3239 747
rect 3876 746 3879 748
rect 3903 746 3913 748
rect 3918 746 3944 748
rect 3956 746 3959 748
rect 3876 736 3879 738
rect 3903 736 3912 738
rect 4385 746 4388 748
rect 4428 746 4446 748
rect 4466 746 4470 748
rect 3917 736 3944 738
rect 3956 736 3959 738
rect 3042 727 3046 728
rect 3018 725 3021 727
rect 3031 725 3046 727
rect 3042 723 3046 725
rect 3042 721 3053 723
rect 3078 721 3081 723
rect 3120 718 3123 720
rect 3133 718 3147 720
rect 3034 713 3053 715
rect 3078 713 3081 715
rect 3145 714 3147 718
rect 3145 712 3155 714
rect 3180 712 3183 714
rect 3120 710 3123 712
rect 3133 710 3142 712
rect 3217 702 3220 704
rect 3230 702 3252 704
rect 3277 702 3280 704
rect 3703 697 3705 700
rect 3872 697 3875 699
rect 3887 697 3901 699
rect 3907 697 3910 699
rect 3927 697 3930 699
rect 3942 697 3956 699
rect 3962 697 3965 699
rect 3018 689 3021 691
rect 3031 689 3045 691
rect 3043 685 3045 689
rect 3742 693 3744 696
rect 3752 693 3754 696
rect 3043 683 3053 685
rect 3078 683 3081 685
rect 3018 681 3021 683
rect 3031 681 3040 683
rect 2935 670 2939 671
rect 2911 668 2914 670
rect 2924 668 2939 670
rect 2935 666 2939 668
rect 3703 671 3705 685
rect 3120 667 3123 669
rect 3133 667 3155 669
rect 3180 667 3183 669
rect 2935 664 2946 666
rect 2971 664 2974 666
rect 3770 687 3772 690
rect 3780 687 3782 690
rect 3703 662 3705 665
rect 3742 660 3744 669
rect 2927 656 2946 658
rect 2971 656 2974 658
rect 3752 659 3754 669
rect 3018 645 3021 647
rect 3031 645 3045 647
rect 3043 641 3045 645
rect 3703 642 3705 645
rect 3043 639 3053 641
rect 3078 639 3081 641
rect 3018 637 3021 639
rect 3031 637 3040 639
rect 2911 632 2914 634
rect 2924 632 2938 634
rect 2936 628 2938 632
rect 2936 626 2946 628
rect 2971 626 2974 628
rect 2911 624 2914 626
rect 2924 624 2933 626
rect 3703 616 3705 630
rect 3742 628 3744 655
rect 3752 628 3754 654
rect 3770 652 3772 663
rect 3770 628 3772 648
rect 3780 641 3782 663
rect 4679 657 4681 660
rect 3780 628 3782 637
rect 4726 638 4728 641
rect 4734 638 4736 641
rect 4764 638 4766 641
rect 4808 638 4810 641
rect 4853 638 4855 641
rect 3742 613 3744 616
rect 3752 613 3754 616
rect 3770 613 3772 616
rect 3780 613 3782 616
rect 3703 607 3705 610
rect 4679 599 4681 617
rect 4891 630 4893 633
rect 4726 606 4728 613
rect 4721 602 4728 606
rect 3018 594 3021 596
rect 3031 594 3053 596
rect 3078 594 3081 596
rect 2911 588 2914 590
rect 2924 588 2938 590
rect 4542 591 4545 593
rect 4595 591 4618 593
rect 2936 584 2938 588
rect 2936 582 2946 584
rect 2971 582 2974 584
rect 2911 580 2914 582
rect 2924 580 2933 582
rect 4722 591 4724 602
rect 4734 594 4736 613
rect 4764 605 4766 613
rect 4808 605 4810 613
rect 4758 603 4766 605
rect 4802 603 4810 605
rect 4758 591 4760 603
rect 4766 591 4768 600
rect 4802 591 4804 603
rect 4810 591 4812 600
rect 4853 591 4855 613
rect 4891 592 4893 610
rect 4679 575 4681 579
rect 4722 578 4724 581
rect 4758 578 4760 581
rect 4766 578 4768 581
rect 4802 578 4804 581
rect 4810 578 4812 581
rect 4853 578 4855 581
rect 4891 578 4893 582
rect 3710 572 3712 575
rect 3749 568 3751 571
rect 3759 568 3761 571
rect 3710 546 3712 560
rect 3777 562 3779 565
rect 3787 562 3789 565
rect 2911 537 2914 539
rect 2924 537 2946 539
rect 2971 537 2974 539
rect 3710 537 3712 540
rect 3749 535 3751 544
rect 3759 534 3761 544
rect 4346 556 4349 558
rect 4399 556 4422 558
rect 4172 552 4175 554
rect 4225 552 4248 554
rect 3710 517 3712 520
rect 3710 491 3712 505
rect 3749 503 3751 530
rect 3759 503 3761 529
rect 3777 527 3779 538
rect 3777 503 3779 523
rect 3787 516 3789 538
rect 3998 529 4001 531
rect 4051 529 4074 531
rect 3787 503 3789 512
rect 4509 506 4521 508
rect 4621 506 4624 508
rect 4321 498 4333 500
rect 4433 498 4436 500
rect 3749 488 3751 491
rect 3759 488 3761 491
rect 3777 488 3779 491
rect 3787 488 3789 491
rect 4140 488 4152 490
rect 4252 488 4255 490
rect 3710 482 3712 485
rect 3972 480 3984 482
rect 4084 480 4087 482
rect 4511 397 4523 399
rect 4623 397 4626 399
rect 4319 387 4331 389
rect 4431 387 4434 389
rect 4139 377 4151 379
rect 4251 377 4254 379
rect 3936 369 3938 372
rect 3732 347 3734 350
rect 3743 347 3745 350
rect 3774 340 3776 344
rect 3732 298 3734 327
rect 3743 298 3745 327
rect 3774 306 3776 320
rect 3774 293 3776 296
rect 3732 275 3734 278
rect 3743 275 3745 278
rect 3971 366 3983 368
rect 4083 366 4086 368
rect 3936 257 3938 269
rect 4013 268 4016 270
rect 4116 268 4128 270
rect 3732 238 3734 241
rect 3743 238 3745 241
rect 4070 237 4073 239
rect 4113 237 4131 239
rect 4151 237 4155 239
rect 3774 231 3776 235
rect 3732 189 3734 218
rect 3743 189 3745 218
rect 3774 197 3776 211
rect 3879 208 3882 210
rect 3907 208 3929 210
rect 3939 208 3942 210
rect 3774 184 3776 187
rect 3732 166 3734 169
rect 3743 166 3745 169
rect 3920 165 3929 167
rect 3939 165 3942 167
rect 3879 163 3882 165
rect 3907 163 3917 165
rect 3915 159 3917 163
rect 3915 157 3929 159
rect 3939 157 3942 159
rect 3733 119 3735 122
rect 3744 119 3746 122
rect 3920 121 3929 123
rect 3939 121 3942 123
rect 3879 119 3882 121
rect 3907 119 3917 121
rect 3775 112 3777 116
rect 3915 115 3917 119
rect 3915 113 3929 115
rect 3939 113 3942 115
rect 3733 70 3735 99
rect 3744 70 3746 99
rect 3775 78 3777 92
rect 3879 89 3882 91
rect 3907 89 3926 91
rect 3879 81 3882 83
rect 3907 81 3918 83
rect 3914 79 3918 81
rect 3914 77 3929 79
rect 3939 77 3942 79
rect 3914 76 3918 77
rect 3775 65 3777 68
rect 3733 47 3735 50
rect 3744 47 3746 50
rect 3737 11 3739 14
rect 3748 11 3750 14
rect 3779 4 3781 8
rect 3737 -38 3739 -9
rect 3748 -38 3750 -9
rect 3779 -30 3781 -16
rect 3779 -43 3781 -40
rect 3737 -61 3739 -58
rect 3748 -61 3750 -58
<< polycontact >>
rect 4155 1169 4160 1173
rect 3642 1134 3646 1138
rect 4161 1132 4165 1136
rect 3634 1121 3638 1125
rect 4160 1117 4165 1122
rect 3642 1110 3646 1114
rect 3634 1097 3639 1102
rect 4342 1100 4347 1104
rect 3634 1083 3638 1087
rect 4161 1088 4165 1092
rect 4160 1073 4165 1078
rect 4519 1077 4524 1081
rect 3543 1062 3547 1066
rect 4153 1061 4157 1065
rect 4348 1063 4352 1067
rect 3535 1049 3539 1053
rect 3634 1053 3639 1058
rect 4161 1050 4165 1054
rect 3543 1038 3547 1042
rect 3634 1039 3638 1043
rect 4347 1048 4352 1053
rect 4153 1037 4157 1041
rect 4525 1040 4529 1044
rect 3535 1025 3540 1030
rect 4524 1025 4529 1030
rect 3535 1011 3539 1015
rect 4348 1019 4352 1023
rect 3639 1002 3644 1006
rect 4347 1004 4352 1009
rect 4340 992 4344 996
rect 4525 996 4529 1000
rect 3535 981 3540 986
rect 4348 981 4352 985
rect 4524 981 4529 986
rect 3447 974 3451 978
rect 3535 967 3539 971
rect 3439 961 3443 965
rect 3447 950 3451 954
rect 3695 950 3699 954
rect 3439 937 3444 942
rect 4340 968 4344 972
rect 4517 969 4521 973
rect 3345 933 3349 937
rect 3540 930 3545 934
rect 3943 960 3948 964
rect 4122 962 4126 966
rect 4525 958 4529 962
rect 4111 951 4115 955
rect 4517 945 4521 949
rect 3337 920 3341 924
rect 3439 923 3443 927
rect 3345 909 3349 913
rect 3337 896 3342 901
rect 3439 893 3444 898
rect 3695 895 3699 899
rect 3764 924 3768 928
rect 3949 923 3953 927
rect 3775 913 3779 917
rect 4291 918 4295 922
rect 3948 908 3953 913
rect 4280 907 4284 911
rect 3337 882 3341 886
rect 3439 879 3443 883
rect 3949 879 3953 883
rect 4085 882 4089 886
rect 4140 882 4144 886
rect 4474 888 4478 892
rect 4463 877 4467 881
rect 3948 864 3953 869
rect 3337 852 3342 857
rect 3941 852 3945 856
rect 3241 836 3245 840
rect 3337 838 3341 842
rect 3444 842 3449 846
rect 3949 841 3953 845
rect 3233 823 3237 827
rect 3696 818 3700 822
rect 3241 812 3245 816
rect 4254 838 4258 842
rect 4309 838 4313 842
rect 3144 801 3148 805
rect 3233 799 3238 804
rect 3342 801 3347 805
rect 3941 828 3945 832
rect 4437 808 4441 812
rect 4492 808 4496 812
rect 3136 788 3140 792
rect 3233 785 3237 789
rect 3144 777 3148 781
rect 3136 764 3141 769
rect 3696 763 3700 767
rect 3765 792 3769 796
rect 3776 781 3780 785
rect 3931 773 3935 777
rect 3233 755 3238 760
rect 3136 750 3140 754
rect 3920 762 3924 766
rect 3233 741 3237 745
rect 3042 728 3046 732
rect 3136 720 3141 725
rect 3034 715 3038 719
rect 3042 704 3046 708
rect 3136 706 3140 710
rect 3238 704 3243 708
rect 3034 691 3039 696
rect 3034 677 3038 681
rect 2935 671 2939 675
rect 3699 674 3703 678
rect 3141 669 3146 673
rect 2927 658 2931 662
rect 3894 693 3898 697
rect 3949 693 3953 697
rect 2935 647 2939 651
rect 3034 647 3039 652
rect 2927 634 2932 639
rect 3034 633 3038 637
rect 2927 620 2931 624
rect 3699 619 3703 623
rect 3768 648 3772 652
rect 3779 637 3783 641
rect 3039 596 3044 600
rect 4674 602 4679 607
rect 4717 602 4721 606
rect 2927 590 2932 595
rect 2927 576 2931 580
rect 4730 594 4734 598
rect 4741 602 4745 606
rect 4753 594 4758 599
rect 4768 594 4772 598
rect 4797 594 4802 599
rect 4849 599 4853 604
rect 4812 594 4816 598
rect 3706 549 3710 553
rect 2932 539 2937 543
rect 3706 494 3710 498
rect 3775 523 3779 527
rect 3786 512 3790 516
rect 3728 301 3732 305
rect 3739 308 3743 312
rect 3770 309 3774 313
rect 3728 192 3732 196
rect 3739 199 3743 203
rect 3770 200 3774 204
rect 3916 204 3921 208
rect 3922 167 3926 171
rect 3921 152 3926 157
rect 3922 123 3926 127
rect 3729 73 3733 77
rect 3740 80 3744 84
rect 3921 108 3926 113
rect 3914 96 3918 100
rect 3771 81 3775 85
rect 3922 85 3926 89
rect 3914 72 3918 76
rect 3733 -35 3737 -31
rect 3744 -28 3748 -24
rect 3775 -27 3779 -23
<< metal1 >>
rect 4156 1220 4160 1225
rect 4146 1216 4164 1220
rect 4113 1208 4126 1212
rect 4174 1208 4184 1212
rect 4116 1207 4120 1208
rect 4116 1202 4120 1203
rect 4111 1172 4115 1188
rect 4156 1180 4161 1195
rect 4146 1176 4168 1180
rect 4111 1168 4121 1172
rect 4183 1172 4187 1180
rect 3612 1138 3616 1139
rect 3612 1134 3621 1138
rect 3642 1138 3646 1145
rect 3684 1134 3688 1140
rect 3612 1102 3616 1134
rect 3621 1118 3631 1126
rect 3634 1125 3638 1134
rect 3678 1130 3688 1134
rect 3621 1114 3653 1118
rect 3637 1105 3639 1110
rect 3634 1102 3639 1105
rect 3642 1109 3646 1110
rect 3612 1098 3621 1102
rect 3513 1066 3517 1067
rect 3513 1062 3522 1066
rect 3543 1066 3547 1073
rect 3585 1062 3589 1068
rect 3513 1030 3517 1062
rect 3522 1046 3532 1054
rect 3535 1053 3539 1062
rect 3579 1058 3589 1062
rect 3522 1042 3554 1046
rect 3538 1033 3540 1038
rect 3535 1030 3540 1033
rect 3543 1037 3547 1038
rect 3513 1026 3522 1030
rect 3513 986 3517 1026
rect 3585 1024 3589 1058
rect 3579 1020 3589 1024
rect 3522 1002 3532 1010
rect 3535 1010 3539 1011
rect 3554 1002 3579 1012
rect 3522 999 3579 1002
rect 3540 994 3545 999
rect 3535 990 3545 994
rect 3535 986 3540 990
rect 3417 978 3421 979
rect 3417 974 3426 978
rect 3447 978 3451 985
rect 3513 982 3522 986
rect 3489 974 3493 980
rect 3315 937 3319 938
rect 3315 933 3324 937
rect 3345 937 3349 944
rect 3417 942 3421 974
rect 3426 958 3436 966
rect 3439 965 3443 974
rect 3483 970 3493 974
rect 3426 954 3458 958
rect 3442 945 3444 950
rect 3439 942 3444 945
rect 3447 949 3451 950
rect 3387 933 3391 939
rect 3315 901 3319 933
rect 3324 917 3334 925
rect 3337 924 3341 933
rect 3381 929 3391 933
rect 3324 913 3356 917
rect 3340 904 3342 909
rect 3337 901 3342 904
rect 3345 908 3349 909
rect 3315 897 3324 901
rect 3315 857 3319 897
rect 3387 895 3391 929
rect 3381 891 3391 895
rect 3324 873 3334 881
rect 3337 881 3341 882
rect 3356 873 3381 883
rect 3324 870 3381 873
rect 3342 865 3347 870
rect 3337 861 3347 865
rect 3337 857 3342 861
rect 3315 853 3324 857
rect 3211 840 3215 841
rect 3211 836 3220 840
rect 3241 840 3245 847
rect 3283 836 3287 842
rect 3114 805 3118 806
rect 3114 801 3123 805
rect 3144 805 3148 812
rect 3186 801 3190 807
rect 3114 769 3118 801
rect 3123 785 3133 793
rect 3136 792 3140 801
rect 3180 797 3190 801
rect 3123 781 3155 785
rect 3139 772 3141 777
rect 3136 769 3141 772
rect 3144 776 3148 777
rect 3114 765 3123 769
rect 3012 732 3016 733
rect 3012 728 3021 732
rect 3042 732 3046 739
rect 3084 728 3088 734
rect 3012 696 3016 728
rect 3021 712 3031 720
rect 3034 719 3038 728
rect 3078 724 3088 728
rect 3021 708 3053 712
rect 3037 699 3039 704
rect 3034 696 3039 699
rect 3042 703 3046 704
rect 3012 692 3021 696
rect 2905 675 2909 676
rect 2905 671 2914 675
rect 2935 675 2939 682
rect 2977 671 2981 677
rect 2905 639 2909 671
rect 2914 655 2924 663
rect 2927 662 2931 671
rect 2971 667 2981 671
rect 2914 651 2946 655
rect 2930 642 2932 647
rect 2927 639 2932 642
rect 2935 646 2939 647
rect 2905 635 2914 639
rect 2905 595 2909 635
rect 2977 633 2981 667
rect 2971 629 2981 633
rect 2914 611 2924 619
rect 2927 619 2931 620
rect 2946 611 2971 621
rect 2914 608 2971 611
rect 2932 603 2937 608
rect 2927 599 2937 603
rect 2927 595 2932 599
rect 2905 591 2914 595
rect 2905 544 2909 591
rect 2977 589 2981 629
rect 3012 652 3016 692
rect 3084 690 3088 724
rect 3078 686 3088 690
rect 3021 668 3031 676
rect 3034 676 3038 677
rect 3053 668 3078 678
rect 3021 665 3078 668
rect 3039 660 3044 665
rect 3034 656 3044 660
rect 3034 652 3039 656
rect 3012 648 3021 652
rect 3012 601 3016 648
rect 3084 646 3088 686
rect 3114 725 3118 765
rect 3186 763 3190 797
rect 3180 759 3190 763
rect 3123 741 3133 749
rect 3136 749 3140 750
rect 3155 741 3180 751
rect 3123 738 3180 741
rect 3141 733 3146 738
rect 3136 729 3146 733
rect 3136 725 3141 729
rect 3114 721 3123 725
rect 3114 674 3118 721
rect 3186 719 3190 759
rect 3180 715 3190 719
rect 3123 697 3133 705
rect 3136 705 3140 706
rect 3155 697 3180 707
rect 3123 694 3180 697
rect 3114 670 3123 674
rect 3141 673 3146 694
rect 3186 674 3190 715
rect 3211 804 3215 836
rect 3220 820 3230 828
rect 3233 827 3237 836
rect 3277 832 3287 836
rect 3220 816 3252 820
rect 3236 807 3238 812
rect 3233 804 3238 807
rect 3241 811 3245 812
rect 3211 800 3220 804
rect 3211 760 3215 800
rect 3283 798 3287 832
rect 3277 794 3287 798
rect 3315 806 3319 853
rect 3387 851 3391 891
rect 3381 847 3391 851
rect 3324 829 3334 837
rect 3337 837 3341 838
rect 3356 829 3381 839
rect 3324 826 3381 829
rect 3315 802 3324 806
rect 3342 805 3347 826
rect 3387 806 3391 847
rect 3417 938 3426 942
rect 3417 898 3421 938
rect 3489 936 3493 970
rect 3483 932 3493 936
rect 3426 914 3436 922
rect 3439 922 3443 923
rect 3458 914 3483 924
rect 3426 911 3483 914
rect 3444 906 3449 911
rect 3439 902 3449 906
rect 3439 898 3444 902
rect 3417 894 3426 898
rect 3417 847 3421 894
rect 3489 892 3493 932
rect 3513 935 3517 982
rect 3585 980 3589 1020
rect 3612 1058 3616 1098
rect 3684 1096 3688 1130
rect 3678 1092 3688 1096
rect 3621 1074 3631 1082
rect 3634 1082 3638 1083
rect 3653 1074 3678 1084
rect 3621 1071 3678 1074
rect 3639 1066 3644 1071
rect 3634 1062 3644 1066
rect 3634 1058 3639 1062
rect 3612 1054 3621 1058
rect 3612 1007 3616 1054
rect 3684 1052 3688 1092
rect 3678 1048 3688 1052
rect 3621 1030 3631 1038
rect 3634 1038 3638 1039
rect 3653 1030 3678 1040
rect 3621 1027 3678 1030
rect 3612 1003 3621 1007
rect 3639 1006 3644 1027
rect 3684 1007 3688 1048
rect 4111 1127 4115 1168
rect 4155 1148 4160 1169
rect 4178 1168 4187 1172
rect 4121 1145 4178 1148
rect 4121 1135 4146 1145
rect 4161 1136 4165 1137
rect 4168 1137 4178 1145
rect 4111 1123 4121 1127
rect 4111 1083 4115 1123
rect 4183 1121 4187 1168
rect 4343 1159 4347 1164
rect 4333 1155 4351 1159
rect 4300 1147 4313 1151
rect 4361 1147 4371 1151
rect 4303 1146 4307 1147
rect 4303 1141 4307 1142
rect 4178 1117 4187 1121
rect 4520 1135 4524 1140
rect 4160 1113 4165 1117
rect 4155 1109 4165 1113
rect 4155 1104 4160 1109
rect 4121 1101 4178 1104
rect 4121 1091 4146 1101
rect 4161 1092 4165 1093
rect 4168 1093 4178 1101
rect 4111 1079 4121 1083
rect 4111 1045 4115 1079
rect 4183 1077 4187 1117
rect 4178 1073 4187 1077
rect 4153 1065 4157 1066
rect 4160 1070 4165 1073
rect 4160 1065 4162 1070
rect 4146 1057 4178 1061
rect 4111 1041 4121 1045
rect 4161 1041 4165 1050
rect 4168 1049 4178 1057
rect 4183 1041 4187 1073
rect 4111 1035 4115 1041
rect 3944 1020 3948 1025
rect 3934 1016 3952 1020
rect 3901 1008 3914 1012
rect 3962 1008 3972 1012
rect 3612 995 3616 1003
rect 3678 1003 3688 1007
rect 3631 995 3653 999
rect 3638 993 3643 995
rect 3684 987 3688 1003
rect 3904 1007 3908 1008
rect 3904 1002 3908 1003
rect 3638 986 3643 987
rect 3579 976 3589 980
rect 3693 979 3721 982
rect 3522 958 3532 966
rect 3535 966 3539 967
rect 3554 958 3579 968
rect 3522 955 3579 958
rect 3513 931 3522 935
rect 3540 934 3545 955
rect 3585 935 3589 976
rect 3694 973 3697 979
rect 3718 978 3721 979
rect 3718 975 3789 978
rect 3643 949 3680 952
rect 3685 950 3695 953
rect 3703 953 3706 961
rect 3733 969 3736 975
rect 3752 969 3755 975
rect 3703 950 3724 953
rect 3703 947 3706 950
rect 3694 937 3697 941
rect 3513 923 3517 931
rect 3579 931 3589 935
rect 3688 935 3712 937
rect 3688 934 3706 935
rect 3532 923 3554 927
rect 3539 920 3544 923
rect 3585 915 3589 931
rect 3711 934 3712 935
rect 3721 927 3724 950
rect 3762 969 3782 972
rect 3762 963 3765 969
rect 3779 963 3782 969
rect 3899 963 3903 979
rect 3944 971 3949 995
rect 4153 985 4157 1037
rect 4178 1037 4187 1041
rect 4183 1036 4187 1037
rect 4298 1103 4302 1119
rect 4343 1111 4348 1134
rect 4510 1131 4528 1135
rect 4477 1123 4490 1127
rect 4538 1123 4548 1127
rect 4480 1122 4484 1123
rect 4480 1117 4484 1118
rect 4333 1107 4355 1111
rect 4298 1099 4308 1103
rect 4370 1103 4374 1111
rect 4298 1058 4302 1099
rect 4342 1079 4347 1100
rect 4365 1099 4374 1103
rect 4308 1076 4365 1079
rect 4308 1066 4333 1076
rect 4348 1067 4352 1068
rect 4355 1068 4365 1076
rect 4298 1054 4308 1058
rect 4121 981 4157 985
rect 4298 1014 4302 1054
rect 4370 1052 4374 1099
rect 4365 1048 4374 1052
rect 4347 1044 4352 1048
rect 4342 1040 4352 1044
rect 4342 1035 4347 1040
rect 4308 1032 4365 1035
rect 4308 1022 4333 1032
rect 4348 1023 4352 1024
rect 4355 1024 4365 1032
rect 4298 1010 4308 1014
rect 3934 967 3956 971
rect 3743 942 3746 945
rect 3743 939 3761 942
rect 3899 959 3909 963
rect 3971 963 3975 971
rect 3771 932 3774 939
rect 3771 929 3788 932
rect 3693 926 3712 927
rect 3688 924 3712 926
rect 3721 924 3764 927
rect 3694 918 3697 924
rect 3785 918 3788 929
rect 3899 918 3903 959
rect 3943 939 3948 960
rect 3966 959 3975 963
rect 3909 936 3966 939
rect 3909 926 3934 936
rect 3949 927 3953 928
rect 3956 928 3966 936
rect 3750 913 3775 916
rect 3785 914 3798 918
rect 3750 911 3753 913
rect 3544 895 3680 898
rect 3685 895 3695 898
rect 3703 898 3706 906
rect 3715 908 3753 911
rect 3785 910 3788 914
rect 3715 898 3718 908
rect 3756 907 3788 910
rect 3756 904 3759 907
rect 3703 895 3718 898
rect 3703 892 3706 895
rect 3483 888 3493 892
rect 3426 870 3436 878
rect 3439 878 3443 879
rect 3458 870 3483 880
rect 3426 867 3483 870
rect 3417 843 3426 847
rect 3444 846 3449 867
rect 3489 847 3493 888
rect 3755 901 3761 904
rect 3694 882 3697 886
rect 3715 885 3720 888
rect 3733 888 3736 892
rect 3780 888 3783 892
rect 3725 885 3789 888
rect 3715 882 3718 885
rect 3688 879 3718 882
rect 3794 879 3798 914
rect 3899 914 3909 918
rect 3899 874 3903 914
rect 3971 912 3975 959
rect 3966 908 3975 912
rect 4061 942 4064 976
rect 4121 975 4125 981
rect 4298 976 4302 1010
rect 4370 1008 4374 1048
rect 4365 1004 4374 1008
rect 4340 996 4344 997
rect 4347 1001 4352 1004
rect 4347 996 4349 1001
rect 4333 988 4365 992
rect 4107 972 4132 975
rect 4067 966 4076 969
rect 4067 952 4070 966
rect 4107 961 4110 972
rect 4100 958 4110 961
rect 4067 949 4076 952
rect 4061 939 4070 942
rect 4061 923 4064 939
rect 4097 933 4100 948
rect 4094 930 4100 933
rect 4061 920 4070 923
rect 4061 908 4064 920
rect 4112 911 4115 951
rect 4123 940 4126 962
rect 4129 946 4132 972
rect 4151 970 4154 976
rect 4147 967 4154 970
rect 4135 946 4138 948
rect 4129 943 4138 946
rect 4135 942 4138 943
rect 4123 937 4131 940
rect 3948 904 3953 908
rect 3943 900 3953 904
rect 3943 895 3948 900
rect 3909 892 3966 895
rect 3909 882 3934 892
rect 3949 883 3953 884
rect 3956 884 3966 892
rect 3899 870 3909 874
rect 3694 847 3722 850
rect 3417 835 3421 843
rect 3483 843 3493 847
rect 3436 835 3458 839
rect 3443 832 3448 835
rect 3489 827 3493 843
rect 3695 841 3698 847
rect 3719 846 3722 847
rect 3719 843 3790 846
rect 3448 817 3681 820
rect 3686 818 3696 821
rect 3704 821 3707 829
rect 3734 837 3737 843
rect 3753 837 3756 843
rect 3704 818 3725 821
rect 3704 815 3707 818
rect 3315 794 3319 802
rect 3381 802 3391 806
rect 3695 805 3698 809
rect 3689 803 3713 805
rect 3689 802 3707 803
rect 3334 794 3356 798
rect 3220 776 3230 784
rect 3233 784 3237 785
rect 3252 776 3277 786
rect 3220 773 3277 776
rect 3238 768 3243 773
rect 3233 764 3243 768
rect 3233 760 3238 764
rect 3211 756 3220 760
rect 3211 709 3215 756
rect 3283 754 3287 794
rect 3341 791 3346 794
rect 3387 786 3391 802
rect 3712 802 3713 803
rect 3722 795 3725 818
rect 3763 837 3783 840
rect 3763 831 3766 837
rect 3780 831 3783 837
rect 3899 836 3903 870
rect 3971 868 3975 908
rect 4057 905 4064 908
rect 4086 908 4115 911
rect 4057 884 4060 905
rect 4086 893 4089 908
rect 4128 905 4131 937
rect 4151 923 4154 967
rect 4298 972 4308 976
rect 4348 972 4352 981
rect 4355 980 4365 988
rect 4370 972 4374 1004
rect 4298 966 4302 972
rect 4340 941 4344 968
rect 4365 968 4374 972
rect 4370 967 4374 968
rect 4475 1080 4479 1096
rect 4520 1088 4525 1110
rect 4510 1084 4532 1088
rect 4475 1076 4485 1080
rect 4547 1080 4551 1088
rect 4475 1035 4479 1076
rect 4519 1056 4524 1077
rect 4542 1076 4551 1080
rect 4485 1053 4542 1056
rect 4485 1043 4510 1053
rect 4525 1044 4529 1045
rect 4532 1045 4542 1053
rect 4475 1031 4485 1035
rect 4475 991 4479 1031
rect 4547 1029 4551 1076
rect 4542 1025 4551 1029
rect 4524 1021 4529 1025
rect 4519 1017 4529 1021
rect 4519 1012 4524 1017
rect 4485 1009 4542 1012
rect 4485 999 4510 1009
rect 4525 1000 4529 1001
rect 4532 1001 4542 1009
rect 4475 987 4485 991
rect 4475 953 4479 987
rect 4547 985 4551 1025
rect 4542 981 4551 985
rect 4517 973 4521 974
rect 4524 978 4529 981
rect 4524 973 4526 978
rect 4510 965 4542 969
rect 4475 949 4485 953
rect 4525 949 4529 958
rect 4532 957 4542 965
rect 4547 949 4551 981
rect 4475 943 4479 949
rect 4290 937 4344 941
rect 4147 920 4154 923
rect 4151 912 4154 920
rect 4151 905 4154 907
rect 4128 902 4144 905
rect 4151 902 4160 905
rect 4102 898 4105 899
rect 4102 893 4104 898
rect 4078 890 4092 893
rect 4057 881 4066 884
rect 4057 880 4060 881
rect 3966 864 3975 868
rect 4086 872 4089 882
rect 4102 884 4105 893
rect 4098 881 4105 884
rect 4102 875 4105 881
rect 4112 884 4115 899
rect 4141 893 4144 902
rect 4133 890 4147 893
rect 4112 881 4121 884
rect 4112 880 4115 881
rect 4113 875 4115 880
rect 4141 872 4144 882
rect 4157 884 4160 902
rect 4153 881 4160 884
rect 4157 875 4160 881
rect 4230 898 4233 932
rect 4290 931 4294 937
rect 4276 928 4301 931
rect 4236 922 4245 925
rect 4236 908 4239 922
rect 4276 917 4279 928
rect 4269 914 4279 917
rect 4236 905 4245 908
rect 4230 895 4239 898
rect 4230 879 4233 895
rect 4266 889 4269 904
rect 4263 886 4269 889
rect 4230 876 4239 879
rect 3941 856 3945 857
rect 3948 861 3953 864
rect 3948 856 3950 861
rect 3934 848 3966 852
rect 3899 832 3909 836
rect 3949 832 3953 841
rect 3956 840 3966 848
rect 3971 832 3975 864
rect 3744 810 3747 813
rect 3744 807 3762 810
rect 3899 826 3903 832
rect 3772 800 3775 807
rect 3772 797 3789 800
rect 3694 794 3713 795
rect 3689 792 3713 794
rect 3722 792 3765 795
rect 3695 786 3698 792
rect 3786 786 3789 797
rect 3941 796 3945 828
rect 3966 828 3975 832
rect 3971 827 3975 828
rect 3930 792 3945 796
rect 4022 795 4026 811
rect 4087 803 4090 867
rect 4141 844 4144 867
rect 4230 864 4233 876
rect 4281 867 4284 907
rect 4292 896 4295 918
rect 4298 902 4301 928
rect 4320 926 4323 932
rect 4316 923 4323 926
rect 4304 902 4307 904
rect 4298 899 4307 902
rect 4304 898 4307 899
rect 4292 893 4300 896
rect 4226 861 4233 864
rect 4255 864 4284 867
rect 4140 841 4145 844
rect 4226 840 4229 861
rect 4255 849 4258 864
rect 4297 861 4300 893
rect 4320 879 4323 923
rect 4517 911 4521 945
rect 4542 945 4551 949
rect 4547 944 4551 945
rect 4473 907 4521 911
rect 4316 876 4323 879
rect 4320 868 4323 876
rect 4320 861 4323 863
rect 4413 868 4416 902
rect 4473 901 4477 907
rect 4459 898 4484 901
rect 4419 892 4428 895
rect 4419 878 4422 892
rect 4459 887 4462 898
rect 4452 884 4462 887
rect 4419 875 4428 878
rect 4413 865 4422 868
rect 4297 858 4313 861
rect 4320 858 4329 861
rect 4271 854 4274 855
rect 4271 849 4273 854
rect 4247 846 4261 849
rect 4226 837 4235 840
rect 4226 836 4229 837
rect 4255 828 4258 838
rect 4271 840 4274 849
rect 4267 837 4274 840
rect 4271 831 4274 837
rect 4281 840 4284 855
rect 4310 849 4313 858
rect 4302 846 4316 849
rect 4281 837 4290 840
rect 4281 836 4284 837
rect 4282 831 4284 836
rect 4310 828 4313 838
rect 4326 840 4329 858
rect 4322 837 4329 840
rect 4326 831 4329 837
rect 4413 849 4416 865
rect 4449 859 4452 874
rect 4446 856 4452 859
rect 4413 846 4422 849
rect 4413 834 4416 846
rect 4464 837 4467 877
rect 4475 866 4478 888
rect 4481 872 4484 898
rect 4503 896 4506 902
rect 4499 893 4506 896
rect 4487 872 4490 874
rect 4481 869 4490 872
rect 4487 868 4490 869
rect 4475 863 4483 866
rect 4409 831 4416 834
rect 4438 834 4467 837
rect 4079 799 4097 803
rect 3751 781 3776 784
rect 3786 782 3799 786
rect 3751 779 3754 781
rect 3346 763 3681 766
rect 3686 763 3696 766
rect 3704 766 3707 774
rect 3716 776 3754 779
rect 3786 778 3789 782
rect 3716 766 3719 776
rect 3757 775 3789 778
rect 3757 772 3760 775
rect 3704 763 3719 766
rect 3704 760 3707 763
rect 3277 750 3287 754
rect 3756 769 3762 772
rect 3695 750 3698 754
rect 3716 753 3721 756
rect 3734 756 3737 760
rect 3781 756 3784 760
rect 3726 753 3790 756
rect 3716 750 3719 753
rect 3220 732 3230 740
rect 3233 740 3237 741
rect 3252 732 3277 742
rect 3220 729 3277 732
rect 3211 705 3220 709
rect 3238 708 3243 729
rect 3283 709 3287 750
rect 3689 747 3719 750
rect 3795 749 3799 782
rect 3795 742 3799 744
rect 3870 753 3873 787
rect 3930 786 3934 792
rect 4022 791 4039 795
rect 4126 795 4130 811
rect 4117 791 4130 795
rect 4029 790 4033 791
rect 3916 783 3941 786
rect 3876 777 3885 780
rect 3876 763 3879 777
rect 3916 772 3919 783
rect 3909 769 3919 772
rect 3876 760 3885 763
rect 3870 750 3879 753
rect 3870 734 3873 750
rect 3906 744 3909 759
rect 3903 741 3909 744
rect 3870 731 3879 734
rect 3870 719 3873 731
rect 3921 722 3924 762
rect 3932 751 3935 773
rect 3938 757 3941 783
rect 3960 781 3963 787
rect 4029 785 4033 786
rect 3956 778 3963 781
rect 3944 757 3947 759
rect 3938 754 3947 757
rect 3944 753 3947 754
rect 3932 748 3940 751
rect 3211 697 3215 705
rect 3277 705 3287 709
rect 3866 716 3873 719
rect 3895 719 3924 722
rect 3230 697 3252 701
rect 3237 694 3242 697
rect 3283 689 3287 705
rect 3697 703 3725 706
rect 3698 697 3701 703
rect 3722 702 3725 703
rect 3722 699 3793 702
rect 3114 662 3118 670
rect 3180 670 3190 674
rect 3242 673 3684 676
rect 3689 674 3699 677
rect 3707 677 3710 685
rect 3737 693 3740 699
rect 3756 693 3759 699
rect 3707 674 3728 677
rect 3707 671 3710 674
rect 3133 662 3155 666
rect 3140 659 3145 662
rect 3186 654 3190 670
rect 3698 661 3701 665
rect 3692 659 3716 661
rect 3692 658 3710 659
rect 3715 658 3716 659
rect 3725 651 3728 674
rect 3766 693 3786 696
rect 3766 687 3769 693
rect 3783 687 3786 693
rect 3866 695 3869 716
rect 3895 704 3898 719
rect 3937 716 3940 748
rect 3960 734 3963 778
rect 3956 731 3963 734
rect 3960 723 3963 731
rect 3960 716 3963 718
rect 3937 713 3953 716
rect 3960 713 3969 716
rect 3911 709 3914 710
rect 3911 704 3913 709
rect 3887 701 3901 704
rect 3866 692 3875 695
rect 3866 691 3869 692
rect 3747 666 3750 669
rect 3747 663 3765 666
rect 3895 683 3898 693
rect 3911 695 3914 704
rect 3907 692 3914 695
rect 3911 686 3914 692
rect 3921 695 3924 710
rect 3950 704 3953 713
rect 3942 701 3956 704
rect 3921 692 3930 695
rect 3921 691 3924 692
rect 3922 686 3924 691
rect 3950 683 3953 693
rect 3966 695 3969 713
rect 3962 692 3969 695
rect 3966 686 3969 692
rect 3775 656 3778 663
rect 3775 653 3792 656
rect 3697 650 3716 651
rect 3692 648 3716 650
rect 3725 648 3768 651
rect 3078 642 3088 646
rect 3021 624 3031 632
rect 3034 632 3038 633
rect 3053 624 3078 634
rect 3021 621 3078 624
rect 3012 597 3021 601
rect 3039 600 3044 621
rect 3084 601 3088 642
rect 3698 642 3701 648
rect 3789 642 3792 653
rect 3754 637 3779 640
rect 3789 638 3802 642
rect 3754 635 3757 637
rect 3145 619 3684 622
rect 3689 619 3699 622
rect 3707 622 3710 630
rect 3719 632 3757 635
rect 3789 634 3792 638
rect 3719 622 3722 632
rect 3760 631 3792 634
rect 3760 628 3763 631
rect 3707 619 3722 622
rect 3707 616 3710 619
rect 3759 625 3765 628
rect 3698 606 3701 610
rect 3719 609 3724 612
rect 3737 612 3740 616
rect 3784 612 3787 616
rect 3729 609 3793 612
rect 3719 606 3722 609
rect 3692 603 3722 606
rect 3798 603 3802 638
rect 3012 589 3016 597
rect 3078 597 3088 601
rect 3031 589 3053 593
rect 2971 585 2981 589
rect 2914 567 2924 575
rect 2927 575 2931 576
rect 2946 567 2971 577
rect 2914 564 2971 567
rect 2905 540 2914 544
rect 2932 543 2937 564
rect 2977 544 2981 585
rect 3038 586 3043 589
rect 3084 581 3088 597
rect 3704 578 3732 581
rect 3705 572 3708 578
rect 3729 577 3732 578
rect 3729 574 3800 577
rect 3044 548 3691 551
rect 3696 549 3706 552
rect 3714 552 3717 560
rect 3744 568 3747 574
rect 3763 568 3766 574
rect 3714 549 3735 552
rect 3714 546 3717 549
rect 2905 532 2909 540
rect 2971 540 2981 544
rect 2924 532 2946 536
rect 2931 529 2936 532
rect 2977 524 2981 540
rect 3705 536 3708 540
rect 3699 534 3723 536
rect 3699 533 3717 534
rect 3722 533 3723 534
rect 3732 526 3735 549
rect 3773 568 3793 571
rect 3773 562 3776 568
rect 3790 562 3793 568
rect 3754 541 3757 544
rect 3754 538 3772 541
rect 3782 531 3785 538
rect 3896 534 3899 678
rect 3948 610 3953 678
rect 3990 541 3995 542
rect 3990 536 3995 537
rect 3985 535 4001 536
rect 3982 534 4001 535
rect 3896 532 4001 534
rect 3896 531 3985 532
rect 3782 528 3799 531
rect 3704 525 3723 526
rect 3699 523 3723 525
rect 3732 523 3775 526
rect 3705 517 3708 523
rect 3796 517 3799 528
rect 3761 512 3786 515
rect 3796 513 3809 517
rect 3761 510 3764 512
rect 2936 494 3691 497
rect 3696 494 3706 497
rect 3714 497 3717 505
rect 3726 507 3764 510
rect 3796 509 3799 513
rect 3726 497 3729 507
rect 3767 506 3799 509
rect 3767 503 3770 506
rect 3714 494 3729 497
rect 3714 491 3717 494
rect 3766 500 3772 503
rect 3705 481 3708 485
rect 3726 484 3731 487
rect 3744 487 3747 491
rect 3791 487 3794 491
rect 3736 484 3800 487
rect 3726 481 3729 484
rect 3699 478 3729 481
rect 3805 476 3809 513
rect 3727 358 3750 362
rect 3731 356 3750 358
rect 3727 347 3731 352
rect 3746 347 3750 356
rect 3763 351 3787 352
rect 3763 347 3779 351
rect 3783 347 3787 351
rect 3763 345 3787 347
rect 3769 340 3773 345
rect 3738 319 3742 327
rect 3738 315 3750 319
rect 3746 313 3750 315
rect 3777 313 3781 320
rect 2931 308 3038 312
rect 3043 308 3739 312
rect 3746 309 3770 313
rect 3777 309 3800 313
rect 2936 301 3728 305
rect 3746 298 3750 309
rect 3777 306 3781 309
rect 3784 308 3800 309
rect 3769 292 3773 296
rect 3763 291 3788 292
rect 3763 287 3783 291
rect 3763 286 3788 287
rect 3727 274 3731 278
rect 3727 270 3743 274
rect 3898 270 3901 531
rect 3990 518 3995 532
rect 4089 528 4093 759
rect 4189 752 4193 772
rect 4256 760 4259 823
rect 4310 818 4313 823
rect 4409 810 4412 831
rect 4438 819 4441 834
rect 4480 831 4483 863
rect 4503 849 4506 893
rect 4499 846 4506 849
rect 4503 838 4506 846
rect 4503 831 4506 833
rect 4480 828 4496 831
rect 4503 828 4512 831
rect 4454 824 4457 825
rect 4454 819 4456 824
rect 4430 816 4444 819
rect 4409 807 4418 810
rect 4409 806 4412 807
rect 4438 798 4441 808
rect 4454 810 4457 819
rect 4450 807 4457 810
rect 4454 801 4457 807
rect 4464 810 4467 825
rect 4493 819 4496 828
rect 4485 816 4499 819
rect 4464 807 4473 810
rect 4464 806 4467 807
rect 4465 801 4467 806
rect 4493 798 4496 808
rect 4509 810 4512 828
rect 4505 807 4512 810
rect 4509 801 4512 807
rect 4246 756 4264 760
rect 4189 748 4206 752
rect 4293 752 4297 772
rect 4284 748 4297 752
rect 4189 741 4193 748
rect 4196 747 4200 748
rect 4196 742 4200 743
rect 4293 741 4297 748
rect 4371 745 4375 761
rect 4439 753 4442 793
rect 4493 790 4496 793
rect 4493 784 4498 790
rect 4428 749 4446 753
rect 4371 741 4388 745
rect 4475 745 4479 761
rect 4466 741 4479 745
rect 4371 733 4375 741
rect 4378 740 4382 741
rect 4378 735 4382 736
rect 4475 733 4479 741
rect 4256 709 4261 715
rect 4164 564 4169 565
rect 4164 559 4169 560
rect 4155 555 4175 559
rect 4164 541 4169 555
rect 4257 551 4261 709
rect 4438 698 4443 702
rect 4439 683 4442 698
rect 4338 568 4343 569
rect 4338 563 4343 564
rect 4329 559 4349 563
rect 4225 547 4261 551
rect 4051 524 4093 528
rect 4089 487 4093 524
rect 4257 497 4261 547
rect 4338 545 4343 559
rect 4438 555 4442 683
rect 4666 670 4687 674
rect 4674 667 4678 670
rect 4668 663 4669 667
rect 4673 663 4678 667
rect 4674 657 4678 663
rect 4715 644 4868 648
rect 4534 603 4539 604
rect 4628 602 4674 607
rect 4682 606 4686 617
rect 4721 638 4725 644
rect 4759 638 4763 644
rect 4803 638 4807 644
rect 4848 638 4852 644
rect 4886 640 4890 643
rect 4771 613 4784 638
rect 4815 613 4828 638
rect 4880 636 4881 640
rect 4885 636 4890 640
rect 4682 602 4717 606
rect 4534 598 4539 599
rect 4525 594 4545 598
rect 4534 580 4539 594
rect 4628 590 4632 602
rect 4682 599 4686 602
rect 4595 586 4632 590
rect 4399 551 4442 555
rect 4438 505 4442 551
rect 4628 513 4632 586
rect 4721 594 4730 598
rect 4737 591 4741 613
rect 4745 602 4746 606
rect 4781 604 4784 613
rect 4825 604 4828 613
rect 4781 599 4793 604
rect 4825 599 4849 604
rect 4856 603 4860 613
rect 4886 630 4890 636
rect 4745 597 4753 599
rect 4750 594 4753 597
rect 4772 594 4773 598
rect 4781 591 4784 599
rect 4789 594 4797 599
rect 4816 594 4817 598
rect 4825 591 4828 599
rect 4856 598 4869 603
rect 4894 600 4898 610
rect 4856 591 4860 598
rect 4894 596 4903 600
rect 4894 592 4898 596
rect 4729 581 4741 591
rect 4773 581 4784 591
rect 4817 581 4828 591
rect 4674 570 4678 579
rect 4717 576 4721 581
rect 4753 576 4757 581
rect 4797 576 4801 581
rect 4848 576 4852 581
rect 4716 572 4860 576
rect 4886 572 4890 582
rect 4666 566 4683 570
rect 4621 509 4632 513
rect 4433 501 4521 505
rect 4256 495 4333 497
rect 4252 493 4333 495
rect 4252 491 4260 493
rect 4084 483 4152 487
rect 3882 265 3901 270
rect 3931 475 3984 479
rect 3931 369 3935 475
rect 4089 373 4093 483
rect 4256 384 4260 491
rect 4437 394 4441 501
rect 4628 404 4632 509
rect 4623 400 4632 404
rect 4431 390 4441 394
rect 4516 392 4523 396
rect 4251 380 4260 384
rect 4325 382 4331 386
rect 4083 369 4093 373
rect 4145 372 4151 376
rect 3977 361 3983 365
rect 3727 249 3750 253
rect 3731 247 3750 249
rect 3727 238 3731 243
rect 3746 238 3750 247
rect 3882 246 3887 265
rect 3898 262 3901 265
rect 3939 267 3943 269
rect 3978 356 3982 361
rect 4145 356 4149 372
rect 4325 356 4329 382
rect 4516 356 4520 392
rect 3978 352 4520 356
rect 3978 267 3982 352
rect 4116 271 4122 275
rect 3939 263 4016 267
rect 3763 242 3787 243
rect 3763 238 3779 242
rect 3783 238 3787 242
rect 3882 241 3922 246
rect 3763 236 3787 238
rect 3769 231 3773 236
rect 3738 210 3742 218
rect 3738 206 3750 210
rect 3746 204 3750 206
rect 3777 204 3781 211
rect 3872 207 3876 223
rect 3917 215 3922 241
rect 4056 236 4060 245
rect 4113 242 4123 244
rect 4128 242 4131 244
rect 4113 240 4131 242
rect 4056 232 4073 236
rect 4160 236 4164 241
rect 4151 232 4164 236
rect 4056 222 4060 232
rect 4063 231 4067 232
rect 4063 226 4067 227
rect 4160 223 4164 232
rect 3907 211 3929 215
rect 3145 199 3739 203
rect 3746 200 3770 204
rect 3777 200 3813 204
rect 3872 203 3882 207
rect 3944 207 3948 215
rect 3141 192 3237 196
rect 3242 192 3728 196
rect 3746 189 3750 200
rect 3777 197 3781 200
rect 3769 183 3773 187
rect 3763 182 3788 183
rect 3763 178 3783 182
rect 3763 177 3788 178
rect 3727 165 3731 169
rect 3727 161 3743 165
rect 3872 162 3876 203
rect 3916 183 3921 204
rect 3939 203 3948 207
rect 3882 180 3939 183
rect 3882 170 3907 180
rect 3922 171 3926 172
rect 3929 172 3939 180
rect 3872 158 3882 162
rect 3728 130 3751 134
rect 3732 128 3751 130
rect 3728 119 3732 124
rect 3747 119 3751 128
rect 3764 123 3788 124
rect 3764 119 3780 123
rect 3784 119 3788 123
rect 3764 117 3788 119
rect 3872 118 3876 158
rect 3944 156 3948 203
rect 3939 152 3948 156
rect 3921 148 3926 152
rect 3916 144 3926 148
rect 3916 139 3921 144
rect 3882 136 3939 139
rect 3882 126 3907 136
rect 3922 127 3926 128
rect 3929 128 3939 136
rect 3770 112 3774 117
rect 3872 114 3882 118
rect 3739 91 3743 99
rect 3739 87 3751 91
rect 3747 85 3751 87
rect 3778 85 3782 92
rect 3333 80 3443 84
rect 3448 80 3740 84
rect 3747 81 3771 85
rect 3778 81 3825 85
rect 3333 73 3341 77
rect 3346 73 3729 77
rect 3747 70 3751 81
rect 3778 78 3782 81
rect 3872 80 3876 114
rect 3944 112 3948 152
rect 3939 108 3948 112
rect 3914 100 3918 101
rect 3921 105 3926 108
rect 3921 100 3923 105
rect 3907 92 3939 96
rect 3872 76 3882 80
rect 3922 76 3926 85
rect 3929 84 3939 92
rect 3944 76 3948 108
rect 3872 70 3876 76
rect 3770 64 3774 68
rect 3914 65 3918 72
rect 3939 72 3948 76
rect 3944 71 3948 72
rect 3764 63 3789 64
rect 3764 59 3784 63
rect 3764 58 3789 59
rect 3728 46 3732 50
rect 3728 42 3744 46
rect 3732 22 3755 26
rect 3736 20 3755 22
rect 3732 11 3736 16
rect 3751 11 3755 20
rect 3768 15 3792 16
rect 3768 11 3784 15
rect 3788 11 3792 15
rect 3768 9 3792 11
rect 3774 4 3778 9
rect 3743 -17 3747 -9
rect 3743 -21 3755 -17
rect 3751 -23 3755 -21
rect 3782 -23 3786 -16
rect 3537 -28 3638 -24
rect 3643 -28 3744 -24
rect 3751 -27 3775 -23
rect 3782 -27 3839 -23
rect 3537 -35 3538 -31
rect 3545 -35 3733 -31
rect 3751 -38 3755 -27
rect 3782 -30 3786 -27
rect 3774 -44 3778 -40
rect 3768 -45 3793 -44
rect 3768 -49 3788 -45
rect 3768 -50 3793 -49
rect 3732 -62 3736 -58
rect 3732 -66 3748 -62
<< m2contact >>
rect 4156 1195 4161 1202
rect 3634 1134 3639 1139
rect 3632 1105 3637 1110
rect 3642 1104 3647 1109
rect 3535 1062 3540 1067
rect 3533 1033 3538 1038
rect 3543 1032 3548 1037
rect 3535 1005 3540 1010
rect 3439 974 3444 979
rect 3337 933 3342 938
rect 3437 945 3442 950
rect 3447 944 3452 949
rect 3335 904 3340 909
rect 3345 903 3350 908
rect 3337 876 3342 881
rect 3233 836 3238 841
rect 3136 801 3141 806
rect 3134 772 3139 777
rect 3144 771 3149 776
rect 3034 728 3039 733
rect 3032 699 3037 704
rect 3042 698 3047 703
rect 2927 671 2932 676
rect 2925 642 2930 647
rect 2935 641 2940 646
rect 2927 614 2932 619
rect 3034 671 3039 676
rect 3136 744 3141 749
rect 3136 700 3141 705
rect 3231 807 3236 812
rect 3241 806 3246 811
rect 3337 832 3342 837
rect 3439 917 3444 922
rect 3634 1077 3639 1082
rect 3634 1033 3639 1038
rect 4160 1137 4165 1142
rect 4343 1134 4348 1140
rect 4160 1093 4165 1098
rect 4152 1066 4157 1071
rect 4162 1065 4167 1070
rect 3638 987 3643 993
rect 3944 995 3949 1002
rect 3535 961 3540 966
rect 3638 948 3643 953
rect 3680 948 3685 953
rect 3539 914 3544 920
rect 4160 1036 4165 1041
rect 4347 1068 4352 1073
rect 4520 1110 4525 1117
rect 4347 1024 4352 1029
rect 3948 928 3953 933
rect 3539 895 3544 900
rect 3680 894 3685 899
rect 3439 873 3444 878
rect 3794 874 3799 879
rect 4339 997 4344 1002
rect 4349 996 4354 1001
rect 3948 884 3953 889
rect 3443 826 3448 832
rect 3443 817 3448 822
rect 3681 816 3686 821
rect 3233 779 3238 784
rect 3341 785 3346 791
rect 4347 967 4352 972
rect 4524 1045 4529 1050
rect 4524 1001 4529 1006
rect 4516 974 4521 979
rect 4526 973 4531 978
rect 4086 867 4091 872
rect 4140 867 4145 872
rect 3940 857 3945 862
rect 3950 856 3955 861
rect 3948 827 3953 832
rect 4140 836 4145 841
rect 4524 944 4529 949
rect 4255 823 4260 828
rect 4309 823 4314 828
rect 3341 763 3346 768
rect 3681 762 3686 767
rect 3233 735 3238 740
rect 3794 744 3799 749
rect 3237 688 3242 694
rect 3237 673 3242 678
rect 3684 672 3689 677
rect 3140 653 3145 659
rect 4089 759 4094 765
rect 3895 678 3900 683
rect 3949 678 3954 683
rect 3034 627 3039 632
rect 3140 619 3145 624
rect 3684 618 3689 623
rect 3798 598 3803 603
rect 2927 570 2932 575
rect 3038 580 3043 586
rect 3039 547 3044 552
rect 3691 547 3696 552
rect 2931 523 2936 529
rect 3948 605 3953 610
rect 2931 493 2936 498
rect 3691 493 3696 498
rect 3805 471 3810 476
rect 3038 308 3043 313
rect 2931 300 2936 305
rect 3800 308 3805 313
rect 4310 812 4316 818
rect 4438 793 4443 798
rect 4492 793 4497 798
rect 4493 778 4498 784
rect 4256 715 4261 723
rect 4438 702 4443 708
rect 4716 594 4721 599
rect 4746 602 4751 607
rect 4745 592 4750 597
rect 4773 594 4778 599
rect 4817 594 4822 599
rect 3898 257 3903 262
rect 4123 242 4128 247
rect 3140 199 3145 204
rect 3813 200 3818 205
rect 3237 191 3242 196
rect 3921 172 3926 177
rect 3921 128 3926 133
rect 3443 80 3448 85
rect 3825 81 3831 87
rect 3341 72 3346 77
rect 3913 101 3918 106
rect 3923 100 3928 105
rect 3921 71 3926 76
rect 3638 -28 3643 -23
rect 3839 -27 3844 -21
rect 3538 -36 3545 -31
<< pm12contact >>
rect 4156 1208 4161 1213
rect 4343 1147 4348 1152
rect 3944 1008 3949 1013
rect 4520 1123 4525 1128
rect 3736 931 3741 936
rect 3745 930 3750 935
rect 4104 932 4109 937
rect 4103 923 4108 928
rect 4273 888 4278 893
rect 4272 879 4277 884
rect 3737 799 3742 804
rect 3746 798 3751 803
rect 4456 858 4461 863
rect 4455 849 4460 854
rect 4089 791 4094 796
rect 3913 743 3918 748
rect 3912 734 3917 739
rect 3740 655 3745 660
rect 3749 654 3754 659
rect 3747 530 3752 535
rect 3756 529 3761 534
rect 4068 531 4074 537
rect 4256 748 4261 753
rect 4438 741 4443 746
rect 4242 554 4248 560
rect 4416 558 4422 564
rect 4612 593 4618 599
rect 4886 595 4891 600
rect 4509 508 4514 513
rect 4321 500 4326 505
rect 4140 490 4145 495
rect 3972 482 3977 487
rect 4511 399 4516 404
rect 4319 389 4324 394
rect 4139 379 4144 384
rect 3971 368 3976 373
rect 4123 263 4128 268
rect 3931 257 3936 262
rect 4123 232 4128 237
<< metal2 >>
rect 4156 1202 4161 1208
rect 3634 1148 3638 1160
rect 3607 1142 3638 1148
rect 4189 1142 4192 1146
rect 3607 1109 3610 1142
rect 3634 1139 3638 1142
rect 4165 1137 4192 1142
rect 3607 1105 3632 1109
rect 3535 1076 3539 1088
rect 3508 1070 3539 1076
rect 3508 1037 3511 1070
rect 3535 1067 3539 1070
rect 3607 1038 3610 1105
rect 3647 1105 3695 1109
rect 3692 1082 3695 1105
rect 3639 1078 3695 1082
rect 4104 1093 4160 1097
rect 4104 1070 4107 1093
rect 4104 1066 4152 1070
rect 4189 1070 4192 1137
rect 4343 1140 4348 1147
rect 4520 1117 4525 1123
rect 4376 1073 4379 1077
rect 4167 1066 4192 1070
rect 4352 1068 4379 1073
rect 3508 1033 3533 1037
rect 3439 988 3443 1000
rect 3412 982 3443 988
rect 3337 947 3341 959
rect 3310 941 3341 947
rect 3310 908 3313 941
rect 3337 938 3341 941
rect 3412 949 3415 982
rect 3439 979 3443 982
rect 3508 966 3511 1033
rect 3548 1033 3596 1037
rect 3593 1010 3596 1033
rect 3607 1033 3634 1038
rect 4161 1033 4165 1036
rect 4189 1033 4192 1066
rect 3607 1029 3610 1033
rect 4161 1027 4192 1033
rect 4161 1015 4165 1027
rect 4291 1024 4347 1028
rect 3540 1006 3596 1010
rect 3944 1002 3949 1008
rect 4291 1001 4294 1024
rect 4291 997 4339 1001
rect 4376 1001 4379 1068
rect 4553 1050 4556 1054
rect 4529 1045 4556 1050
rect 4354 997 4379 1001
rect 3638 993 3643 995
rect 3508 961 3535 966
rect 3508 957 3511 961
rect 3638 953 3643 987
rect 4348 964 4352 967
rect 4376 964 4379 997
rect 4468 1001 4524 1005
rect 4468 978 4471 1001
rect 4468 974 4516 978
rect 4553 978 4556 1045
rect 4531 974 4556 978
rect 4348 958 4379 964
rect 3412 945 3437 949
rect 3310 904 3335 908
rect 3233 850 3237 862
rect 3206 844 3237 850
rect 3136 815 3140 827
rect 3109 809 3140 815
rect 3109 776 3112 809
rect 3136 806 3140 809
rect 3206 811 3209 844
rect 3233 841 3237 844
rect 3310 837 3313 904
rect 3350 904 3398 908
rect 3395 881 3398 904
rect 3342 877 3398 881
rect 3412 878 3415 945
rect 3452 945 3500 949
rect 3497 922 3500 945
rect 3444 918 3500 922
rect 3539 920 3544 923
rect 3539 900 3544 914
rect 3412 873 3439 878
rect 3412 869 3415 873
rect 3310 832 3337 837
rect 3443 832 3448 835
rect 3310 828 3313 832
rect 3443 822 3448 826
rect 3206 807 3231 811
rect 3109 772 3134 776
rect 3034 742 3038 754
rect 3007 736 3038 742
rect 3007 703 3010 736
rect 3034 733 3038 736
rect 3109 705 3112 772
rect 3149 772 3197 776
rect 3194 749 3197 772
rect 3141 745 3197 749
rect 3206 740 3209 807
rect 3246 807 3294 811
rect 3291 784 3294 807
rect 3238 780 3294 784
rect 3341 791 3346 794
rect 3341 768 3346 785
rect 3206 735 3233 740
rect 3206 731 3209 735
rect 3007 699 3032 703
rect 2927 685 2931 697
rect 2900 679 2931 685
rect 2900 646 2903 679
rect 2927 676 2931 679
rect 2900 642 2925 646
rect 2900 575 2903 642
rect 2940 642 2988 646
rect 2985 619 2988 642
rect 3007 632 3010 699
rect 3047 699 3095 703
rect 3092 676 3095 699
rect 3109 700 3136 705
rect 3109 696 3112 700
rect 3039 672 3095 676
rect 3237 694 3242 697
rect 3237 678 3242 688
rect 3007 627 3034 632
rect 3007 623 3010 627
rect 3140 624 3145 653
rect 2932 615 2988 619
rect 3038 586 3043 587
rect 2900 570 2927 575
rect 2900 566 2903 570
rect 3038 552 3043 580
rect 2931 498 2936 523
rect 2931 305 2936 493
rect 2931 299 2936 300
rect 3038 313 3043 547
rect 3038 299 3043 308
rect 3140 204 3145 619
rect 3141 189 3145 199
rect 3237 196 3242 673
rect 3237 189 3242 191
rect 3341 77 3346 763
rect 3443 85 3448 817
rect 3443 72 3448 80
rect 3539 -31 3544 895
rect 3638 -23 3643 948
rect 3681 942 3684 948
rect 4348 946 4352 958
rect 3681 939 3718 942
rect 3715 936 3718 939
rect 4525 941 4529 944
rect 4553 941 4556 974
rect 3715 933 3736 936
rect 3977 933 3980 937
rect 3745 920 3748 930
rect 3953 928 3980 933
rect 4525 935 4556 941
rect 4109 932 4122 935
rect 3682 917 3748 920
rect 3682 899 3685 917
rect 3892 884 3948 888
rect 3799 874 3854 879
rect 3682 810 3685 816
rect 3682 807 3719 810
rect 3716 804 3719 807
rect 3716 801 3737 804
rect 3746 788 3749 798
rect 3683 785 3749 788
rect 3683 767 3686 785
rect 3799 744 3842 749
rect 3685 666 3688 672
rect 3685 663 3722 666
rect 3719 660 3722 663
rect 3719 657 3740 660
rect 3749 644 3752 654
rect 3686 641 3752 644
rect 3686 623 3689 641
rect 3803 599 3821 603
rect 3692 541 3695 547
rect 3692 538 3729 541
rect 3726 535 3729 538
rect 3726 532 3747 535
rect 3756 519 3759 529
rect 3693 516 3759 519
rect 3693 498 3696 516
rect 3805 435 3810 471
rect 3817 445 3821 599
rect 3837 455 3842 744
rect 3849 470 3854 874
rect 3892 861 3895 884
rect 3892 857 3940 861
rect 3977 861 3980 928
rect 4103 905 4106 923
rect 4097 902 4106 905
rect 4097 871 4100 902
rect 4091 868 4100 871
rect 4119 872 4122 932
rect 4525 923 4529 935
rect 4278 888 4291 891
rect 4119 869 4140 872
rect 4272 861 4275 879
rect 3955 857 3980 861
rect 3949 824 3953 827
rect 3977 824 3980 857
rect 4266 858 4275 861
rect 3949 818 3980 824
rect 3949 806 3953 818
rect 4089 765 4094 791
rect 3918 743 3931 746
rect 3912 716 3915 734
rect 3906 713 3915 716
rect 3906 682 3909 713
rect 3900 679 3909 682
rect 3928 683 3931 743
rect 3928 680 3949 683
rect 3953 605 3985 610
rect 3972 495 3977 605
rect 4068 537 4074 541
rect 4140 505 4145 836
rect 4266 827 4269 858
rect 4260 824 4269 827
rect 4288 828 4291 888
rect 4461 858 4474 861
rect 4455 831 4458 849
rect 4449 828 4458 831
rect 4288 825 4309 828
rect 4316 812 4325 816
rect 4256 723 4261 748
rect 4242 560 4248 564
rect 4321 514 4325 812
rect 4449 797 4452 828
rect 4443 794 4452 797
rect 4471 798 4474 858
rect 4471 795 4492 798
rect 4438 708 4443 741
rect 4493 689 4498 778
rect 4493 684 4514 689
rect 4493 683 4498 684
rect 4416 564 4422 568
rect 4509 526 4514 684
rect 4746 652 4777 655
rect 4612 599 4618 603
rect 4746 607 4750 652
rect 4773 599 4777 652
rect 4695 594 4716 598
rect 4707 570 4713 594
rect 4877 595 4886 600
rect 4746 570 4750 592
rect 4817 570 4822 594
rect 4707 567 4826 570
rect 3962 490 3977 495
rect 3962 470 3967 490
rect 3972 487 3977 490
rect 4131 500 4145 505
rect 3849 465 3967 470
rect 4131 455 4136 500
rect 4140 495 4145 500
rect 4312 510 4325 514
rect 3837 450 4136 455
rect 4312 445 4316 510
rect 4321 509 4325 510
rect 4496 521 4514 526
rect 4321 505 4326 509
rect 3817 441 4316 445
rect 4496 435 4501 521
rect 4509 513 4514 521
rect 3805 430 4501 435
rect 3800 406 4516 411
rect 3800 313 3805 406
rect 4511 404 4516 406
rect 3813 396 4324 401
rect 3813 205 3818 396
rect 4319 394 4324 396
rect 3825 385 4144 391
rect 3825 87 3831 385
rect 4139 384 4144 385
rect 3839 376 3976 381
rect 3839 -21 3844 376
rect 3971 373 3976 376
rect 3903 257 3931 262
rect 4123 257 4128 263
rect 4123 247 4128 252
rect 4123 229 4128 232
rect 3950 177 3953 181
rect 3926 172 3953 177
rect 3865 128 3921 132
rect 3865 105 3869 128
rect 3865 101 3913 105
rect 3950 105 3953 172
rect 3928 101 3953 105
rect 3922 68 3926 71
rect 3950 68 3953 101
rect 3922 62 3953 68
rect 3922 50 3926 62
rect 3638 -35 3643 -28
<< m3contact >>
rect 4068 541 4074 547
rect 4242 564 4248 570
rect 4416 568 4422 574
rect 4612 603 4618 609
rect 4123 252 4128 257
<< m123contact >>
rect 3688 979 3693 984
rect 3688 926 3693 931
rect 3706 930 3711 935
rect 3720 885 3725 890
rect 3689 847 3694 852
rect 3689 794 3694 799
rect 3707 798 3712 803
rect 3721 753 3726 758
rect 3692 703 3697 708
rect 3692 650 3697 655
rect 3710 654 3715 659
rect 3724 609 3729 614
rect 3699 578 3704 583
rect 3699 525 3704 530
rect 3717 529 3722 534
rect 3731 484 3736 489
rect 4055 875 4060 880
rect 4104 893 4109 898
rect 4108 875 4113 880
rect 4149 907 4154 912
rect 3864 686 3869 691
rect 3913 704 3918 709
rect 3917 686 3922 691
rect 3958 718 3963 723
rect 4224 831 4229 836
rect 4273 849 4278 854
rect 4277 831 4282 836
rect 4318 863 4323 868
rect 4407 801 4412 806
rect 4456 819 4461 824
rect 4460 801 4465 806
rect 4501 833 4506 838
<< metal3 >>
rect 3688 931 3691 979
rect 3711 930 3723 933
rect 3720 890 3723 930
rect 4106 907 4149 910
rect 4106 898 4109 907
rect 4060 875 4108 878
rect 4275 863 4318 866
rect 4275 854 4278 863
rect 3689 799 3692 847
rect 4229 831 4277 834
rect 4458 833 4501 836
rect 4458 824 4461 833
rect 4412 801 4460 804
rect 3712 798 3724 801
rect 3721 758 3724 798
rect 3915 718 3958 721
rect 3915 709 3918 718
rect 3692 655 3695 703
rect 3869 686 3917 689
rect 3715 654 3727 657
rect 3724 614 3727 654
rect 4068 634 4618 639
rect 3699 530 3702 578
rect 4068 547 4074 634
rect 4242 570 4248 634
rect 3722 529 3734 532
rect 3731 489 3734 529
rect 4280 257 4285 634
rect 4416 574 4422 634
rect 4612 609 4618 634
rect 4128 252 4285 257
<< labels >>
rlabel metal1 4086 369 4091 373 3 pdr1
rlabel metal2 3971 373 3976 377 3 gen_1
rlabel metal1 3931 372 3935 377 1 prop1_car0
rlabel metal2 3927 257 3931 262 1 carry_0
rlabel metal1 3939 263 3943 268 1 clock_car0
rlabel metal1 4008 263 4013 267 7 clock_car0
rlabel metal2 4123 259 4128 263 7 clock_in
rlabel metal1 4117 271 4122 275 7 gnd!
rlabel metal1 3977 361 3982 365 3 clock_car0
rlabel metal1 4088 483 4092 487 3 pdr1
rlabel metal2 3972 487 3977 491 4 prop_1
rlabel metal1 3978 475 3983 479 3 prop1_car0
rlabel space 3981 532 3986 536 3 vdd!
rlabel m3contact 4068 541 4074 547 6 clock_in
rlabel metal1 4060 524 4065 528 7 pdr1
rlabel metal1 4145 372 4150 376 3 clock_car0
rlabel metal2 4139 384 4144 388 3 gen_2
rlabel metal1 4254 380 4259 384 3 pdr2
rlabel metal1 4255 491 4260 495 3 pdr2
rlabel metal2 4140 495 4145 499 3 prop_2
rlabel metal1 4146 483 4151 487 3 pdr1
rlabel metal1 4155 555 4160 559 3 vdd!
rlabel m3contact 4242 564 4248 570 7 clock_in
rlabel metal1 4235 547 4239 551 7 pdr2
rlabel metal1 4325 382 4330 386 3 clock_car0
rlabel metal2 4319 394 4324 398 3 gen_3
rlabel metal1 4434 390 4439 394 3 pdr3
rlabel metal1 4626 400 4631 404 3 pdr4
rlabel metal2 4511 404 4516 408 3 gen_4
rlabel metal1 4517 392 4522 396 1 clock_car0
rlabel metal1 4436 501 4441 505 3 pdr3
rlabel metal2 4321 505 4326 509 3 prop_3
rlabel metal1 4327 493 4332 497 3 pdr2
rlabel metal1 4624 509 4629 513 3 pdr4
rlabel metal2 4509 513 4514 517 3 prop_4
rlabel metal1 4515 501 4520 505 3 pdr3
rlabel metal1 4329 559 4334 563 3 vdd!
rlabel m3contact 4416 568 4422 574 7 clock_in
rlabel metal1 4409 551 4413 555 7 pdr3
rlabel metal1 4525 594 4530 598 3 vdd!
rlabel m3contact 4612 604 4618 609 7 clock_in
rlabel metal1 4605 586 4609 590 7 pdr4
rlabel metal1 4682 602 4686 607 1 c4
rlabel metal1 4675 670 4680 674 5 vdd!
rlabel metal1 4679 566 4683 570 1 gnd!
rlabel metal1 4725 574 4728 575 1 gnd
rlabel metal1 4731 646 4733 647 5 vdd
rlabel metal2 4712 595 4712 595 1 clk_org
rlabel metal1 4712 604 4712 604 1 c4
rlabel metal1 4867 601 4867 601 7 q_c4
rlabel metal1 4889 639 4889 639 5 vdd!
rlabel metal1 4889 575 4889 575 1 gnd!
rlabel metal2 4879 598 4879 598 1 q_c4
rlabel metal1 4901 597 4901 597 7 iq_c4
rlabel metal1 4160 237 4164 241 7 gnd!
rlabel metal1 4056 233 4060 238 3 vdd!
rlabel metal2 4123 229 4128 232 7 clk_org
rlabel metal1 4123 240 4128 244 7 clock_in
rlabel metal1 3742 23 3742 23 5 vdd
rlabel metal1 3743 -64 3743 -64 1 gnd
rlabel metal1 3775 -46 3775 -46 1 gnd
rlabel metal1 3772 11 3772 11 5 vdd
rlabel metal1 3727 -26 3727 -26 3 q_a1
rlabel metal1 3729 -33 3729 -33 3 q_b1
rlabel metal1 3791 -26 3791 -26 1 gen_1
rlabel metal1 3738 131 3738 131 5 vdd
rlabel metal1 3739 44 3739 44 1 gnd
rlabel metal1 3771 62 3771 62 1 gnd
rlabel metal1 3768 119 3768 119 5 vdd
rlabel metal1 3724 81 3724 81 1 q_a2
rlabel metal1 3724 74 3724 74 1 q_b2
rlabel metal1 3787 83 3787 83 1 gen_2
rlabel metal1 3737 250 3737 250 5 vdd
rlabel metal1 3738 163 3738 163 1 gnd
rlabel metal1 3770 181 3770 181 1 gnd
rlabel metal1 3767 238 3767 238 5 vdd
rlabel metal1 3722 200 3722 200 1 q_b3
rlabel metal1 3724 193 3724 193 1 q_a3
rlabel metal1 3785 202 3785 202 1 gen_3
rlabel metal1 3737 359 3737 359 5 vdd
rlabel metal1 3738 272 3738 272 1 gnd
rlabel metal1 3770 290 3770 290 1 gnd
rlabel metal1 3767 347 3767 347 5 vdd
rlabel metal1 3722 310 3722 310 3 q_a4
rlabel metal1 3722 304 3722 304 3 q_b4
rlabel metal1 3785 311 3785 311 1 gen_4
rlabel metal1 3797 785 3797 785 1 prop_2
rlabel metal1 3679 764 3679 764 3 q_b2
rlabel metal1 3679 819 3679 819 3 q_a2
rlabel metal1 3702 793 3705 795 1 vdd
rlabel metal1 3701 847 3704 849 5 vdd
rlabel metal1 3705 803 3706 805 1 gnd
rlabel metal1 3757 753 3760 755 1 gnd
rlabel metal1 3707 747 3711 750 1 gnd
rlabel metal1 3710 603 3714 606 1 gnd
rlabel metal1 3760 609 3763 611 1 gnd
rlabel metal1 3708 659 3709 661 1 gnd
rlabel metal1 3704 703 3707 705 5 vdd
rlabel metal1 3705 649 3708 651 1 vdd
rlabel metal1 3683 675 3683 675 1 q_a3
rlabel metal1 3683 621 3683 621 1 q_b3
rlabel metal1 3800 640 3800 640 1 prop_3
rlabel metal1 3717 478 3721 481 1 gnd
rlabel metal1 3767 484 3770 486 1 gnd
rlabel metal1 3715 534 3716 536 1 gnd
rlabel metal1 3711 578 3714 580 5 vdd
rlabel metal1 3712 524 3715 526 1 vdd
rlabel metal1 3689 549 3689 549 1 q_a4
rlabel metal1 3689 496 3689 496 1 q_b4
rlabel metal1 3808 515 3808 515 1 prop_4
rlabel metal1 3794 916 3794 916 1 prop_1
rlabel metal1 3678 897 3678 897 1 q_b1
rlabel metal1 3678 951 3678 951 1 q_a1
rlabel metal1 3701 925 3704 927 1 vdd
rlabel metal1 3700 979 3703 981 5 vdd
rlabel metal1 3704 935 3705 937 1 gnd
rlabel metal1 3756 885 3759 887 1 gnd
rlabel metal1 3706 879 3710 882 1 gnd
rlabel metal1 3945 80 3946 83 7 gnd
rlabel metal1 3873 86 3874 88 3 vdd
rlabel metal2 3925 67 3925 67 7 clk_org
rlabel metal1 3916 66 3916 66 7 cin
rlabel metal1 3920 223 3920 223 7 carry_0
rlabel metal1 4441 791 4441 791 7 c3
rlabel metal1 4494 791 4494 791 7 prop_4
rlabel metal1 4475 909 4475 909 7 s4
rlabel metal1 4464 814 4466 817 7 vdd
rlabel metal1 4410 813 4412 816 3 vdd
rlabel metal1 4454 817 4456 818 7 gnd
rlabel metal1 4504 869 4506 872 7 gnd
rlabel metal1 4509 819 4512 823 7 gnd
rlabel metal2 4438 738 4443 741 7 pdr3
rlabel metal1 4438 749 4443 753 7 c3
rlabel metal1 4371 741 4375 745 3 vdd!
rlabel metal1 4475 745 4479 749 7 gnd!
rlabel metal1 4126 800 4130 804 7 gnd!
rlabel metal1 4022 791 4026 795 3 vdd!
rlabel metal1 4089 799 4094 803 7 c1
rlabel metal2 4089 788 4094 791 7 pdr1
rlabel metal1 4293 759 4297 763 7 gnd!
rlabel metal1 4189 748 4193 752 3 vdd!
rlabel metal1 4256 756 4261 760 7 c2
rlabel metal2 4256 745 4261 748 7 pdr2
rlabel metal1 3946 1024 3946 1024 7 iq_s1
rlabel m2contact 3947 1001 3947 1001 7 q_s1
rlabel metal1 3969 1011 3969 1011 7 gnd!
rlabel metal1 3905 1011 3905 1011 3 vdd!
rlabel metal1 3946 978 3946 978 5 q_s1
rlabel metal1 3943 823 3943 823 7 s1
rlabel metal2 3952 823 3952 823 7 clk_org
rlabel metal1 3900 842 3901 844 3 vdd
rlabel metal1 3972 836 3973 839 7 gnd
rlabel metal1 3932 795 3932 795 7 s1
rlabel metal1 3951 676 3951 676 7 prop_1
rlabel metal1 3897 676 3897 676 7 carry_0
rlabel metal1 3921 699 3923 702 7 vdd
rlabel metal1 3867 698 3869 701 3 vdd
rlabel metal1 3911 702 3913 703 7 gnd
rlabel metal1 3961 754 3963 757 7 gnd
rlabel metal1 3966 704 3969 708 7 gnd
rlabel metal1 4158 1223 4158 1223 7 iq_s2
rlabel metal2 4159 1202 4159 1202 7 q_s2
rlabel metal1 4181 1211 4181 1211 7 gnd!
rlabel metal1 4117 1211 4117 1211 3 vdd!
rlabel metal1 4159 1186 4159 1186 7 q_s2
rlabel metal1 4155 1033 4155 1033 7 s2
rlabel metal2 4164 1032 4164 1032 7 clk_org
rlabel metal1 4112 1051 4113 1053 3 vdd
rlabel metal1 4184 1045 4185 1048 7 gnd
rlabel metal1 4124 984 4124 984 5 s2
rlabel metal1 4143 865 4143 865 7 prop_2
rlabel metal1 4089 866 4089 866 7 c1
rlabel metal1 4112 888 4114 891 7 vdd
rlabel metal1 4058 887 4060 890 3 vdd
rlabel metal1 4102 891 4104 892 7 gnd
rlabel metal1 4152 943 4154 946 7 gnd
rlabel metal1 4157 893 4160 897 7 gnd
rlabel metal1 4326 849 4329 853 7 gnd
rlabel metal1 4321 899 4323 902 7 gnd
rlabel metal1 4271 847 4273 848 7 gnd
rlabel metal1 4227 843 4229 846 3 vdd
rlabel metal1 4281 844 4283 847 7 vdd
rlabel metal1 4257 821 4257 821 7 c2
rlabel metal1 4292 940 4292 940 7 s3
rlabel metal1 4312 819 4312 819 7 prop_3
rlabel metal1 4371 976 4372 979 7 gnd
rlabel metal1 4299 982 4300 984 3 vdd
rlabel metal2 4351 963 4351 963 7 clk_org
rlabel metal1 4342 963 4342 963 7 s3
rlabel metal1 4345 1118 4345 1118 7 q_s3
rlabel metal1 4304 1150 4304 1150 3 vdd!
rlabel metal1 4368 1150 4368 1150 7 gnd!
rlabel metal2 4346 1140 4346 1140 7 q_s3
rlabel metal1 4345 1162 4345 1162 7 iq_s3
rlabel metal1 4548 953 4549 956 7 gnd
rlabel metal1 4476 959 4477 961 3 vdd
rlabel metal2 4528 940 4528 940 7 clk_org
rlabel metal1 4519 940 4519 940 7 s4
rlabel metal1 4523 1094 4523 1094 7 q_s4
rlabel metal1 4481 1126 4481 1126 3 vdd!
rlabel metal1 4545 1126 4545 1126 7 gnd!
rlabel metal2 4522 1117 4522 1117 7 q_s4
rlabel metal1 4522 1138 4522 1138 7 iq_s4
rlabel m2contact 2934 525 2934 525 3 q_b4
rlabel metal1 2937 680 2937 680 3 b4
rlabel metal2 2928 680 2928 680 3 clk_org
rlabel metal1 2979 659 2980 661 7 vdd
rlabel metal1 2907 664 2908 667 3 gnd
rlabel metal1 3014 721 3015 724 3 gnd
rlabel metal1 3086 716 3087 718 7 vdd
rlabel metal2 3035 737 3035 737 3 clk_org
rlabel metal1 3045 737 3045 737 3 a4
rlabel m2contact 3040 582 3040 582 3 q_a4
rlabel m2contact 3143 654 3143 654 3 q_b3
rlabel metal1 3146 809 3146 809 3 b3
rlabel metal2 3137 810 3137 810 3 clk_org
rlabel metal1 3188 789 3189 791 7 vdd
rlabel metal1 3116 794 3117 797 3 gnd
rlabel metal1 3213 829 3214 832 3 gnd
rlabel metal1 3285 824 3286 826 7 vdd
rlabel metal2 3234 845 3234 845 3 clk_org
rlabel metal1 3243 845 3243 845 3 a3
rlabel m2contact 3239 691 3239 691 3 q_a3
rlabel metal1 3317 926 3318 929 3 gnd
rlabel metal1 3389 921 3390 923 7 vdd
rlabel metal2 3338 942 3338 942 3 clk_org
rlabel metal1 3347 941 3347 941 3 b2
rlabel m2contact 3343 788 3343 788 3 q_b2
rlabel m2contact 3445 828 3445 828 3 q_a2
rlabel metal1 3449 983 3449 983 3 a2
rlabel metal2 3440 983 3440 983 3 clk_org
rlabel metal1 3491 962 3492 964 7 vdd
rlabel metal1 3419 967 3420 970 3 gnd
rlabel m2contact 3542 916 3542 916 3 q_b1
rlabel metal1 3515 1055 3516 1058 3 gnd
rlabel metal1 3587 1050 3588 1052 7 vdd
rlabel metal2 3536 1071 3536 1071 3 clk_org
rlabel metal1 3545 1071 3545 1071 3 b1
rlabel metal1 3614 1127 3615 1130 3 gnd
rlabel metal1 3686 1122 3687 1124 7 vdd
rlabel metal2 3635 1143 3635 1143 3 clk_org
rlabel metal1 3644 1143 3644 1143 3 a1
rlabel m2contact 3641 988 3641 988 3 q_a1
<< end >>
