magic
tech scmos
timestamp 1731947368
<< nwell >>
rect -263 -624 -239 -562
rect -213 -623 -189 -561
rect -163 -623 -139 -561
rect -116 -623 -92 -561
rect 85 -601 109 -549
rect 163 -762 187 -710
rect 201 -762 225 -710
rect 245 -762 269 -710
rect 283 -762 307 -710
<< ntransistor >>
rect 96 -633 98 -613
rect -318 -778 -316 -678
rect -284 -778 -282 -678
rect -249 -777 -247 -677
rect -214 -778 -212 -678
rect -177 -777 -175 -677
rect -140 -776 -138 -676
rect -104 -776 -102 -676
rect -68 -776 -66 -676
rect -34 -775 -32 -675
rect 5 -774 7 -674
rect 174 -794 176 -774
rect 212 -794 214 -774
rect 256 -794 258 -774
rect 294 -794 296 -774
<< ptransistor >>
rect -252 -618 -250 -568
rect -202 -617 -200 -567
rect -152 -617 -150 -567
rect -105 -617 -103 -567
rect 96 -595 98 -555
rect 174 -756 176 -716
rect 212 -756 214 -716
rect 256 -756 258 -716
rect 294 -756 296 -716
<< ndiffusion >>
rect 95 -633 96 -613
rect 98 -633 99 -613
rect -319 -778 -318 -678
rect -316 -778 -315 -678
rect -285 -778 -284 -678
rect -282 -778 -281 -678
rect -250 -777 -249 -677
rect -247 -777 -246 -677
rect -215 -778 -214 -678
rect -212 -778 -211 -678
rect -178 -777 -177 -677
rect -175 -777 -174 -677
rect -141 -776 -140 -676
rect -138 -776 -137 -676
rect -105 -776 -104 -676
rect -102 -776 -101 -676
rect -69 -776 -68 -676
rect -66 -776 -65 -676
rect -35 -775 -34 -675
rect -32 -775 -31 -675
rect 4 -774 5 -674
rect 7 -774 8 -674
rect 173 -794 174 -774
rect 176 -794 177 -774
rect 211 -794 212 -774
rect 214 -794 215 -774
rect 255 -794 256 -774
rect 258 -794 259 -774
rect 293 -794 294 -774
rect 296 -794 297 -774
<< pdiffusion >>
rect -253 -618 -252 -568
rect -250 -618 -249 -568
rect -203 -617 -202 -567
rect -200 -617 -199 -567
rect -153 -617 -152 -567
rect -150 -617 -149 -567
rect -106 -617 -105 -567
rect -103 -617 -102 -567
rect 95 -595 96 -555
rect 98 -595 99 -555
rect 173 -756 174 -716
rect 176 -756 177 -716
rect 211 -756 212 -716
rect 214 -756 215 -716
rect 255 -756 256 -716
rect 258 -756 259 -716
rect 293 -756 294 -716
rect 296 -756 297 -716
<< ndcontact >>
rect 91 -633 95 -613
rect 99 -633 103 -613
rect -323 -778 -319 -678
rect -315 -778 -311 -678
rect -289 -778 -285 -678
rect -281 -778 -277 -678
rect -254 -777 -250 -677
rect -246 -777 -242 -677
rect -219 -778 -215 -678
rect -211 -778 -207 -678
rect -182 -777 -178 -677
rect -174 -777 -170 -677
rect -145 -776 -141 -676
rect -137 -776 -133 -676
rect -109 -776 -105 -676
rect -101 -776 -97 -676
rect -73 -776 -69 -676
rect -65 -776 -61 -676
rect -39 -775 -35 -675
rect -31 -775 -27 -675
rect 0 -774 4 -674
rect 8 -774 12 -674
rect 169 -794 173 -774
rect 177 -794 181 -774
rect 207 -794 211 -774
rect 215 -794 219 -774
rect 251 -794 255 -774
rect 259 -794 263 -774
rect 289 -794 293 -774
rect 297 -794 301 -774
<< pdcontact >>
rect -257 -618 -253 -568
rect -249 -618 -245 -568
rect -207 -617 -203 -567
rect -199 -617 -195 -567
rect -157 -617 -153 -567
rect -149 -617 -145 -567
rect -110 -617 -106 -567
rect -102 -617 -98 -567
rect 91 -595 95 -555
rect 99 -595 103 -555
rect 169 -756 173 -716
rect 177 -756 181 -716
rect 207 -756 211 -716
rect 215 -756 219 -716
rect 251 -756 255 -716
rect 259 -756 263 -716
rect 289 -756 293 -716
rect 297 -756 301 -716
<< nsubstratencontact >>
rect 86 -549 90 -545
rect -262 -562 -258 -557
rect -212 -561 -208 -556
rect -162 -561 -158 -556
rect -115 -561 -111 -556
rect 164 -710 168 -706
rect 202 -710 206 -706
rect 246 -710 250 -706
rect 284 -710 288 -706
<< polysilicon >>
rect 96 -555 98 -552
rect -252 -568 -250 -565
rect -202 -567 -200 -564
rect -152 -567 -150 -564
rect -105 -567 -103 -564
rect 96 -613 98 -595
rect -252 -641 -250 -618
rect -202 -640 -200 -617
rect -152 -640 -150 -617
rect -105 -640 -103 -617
rect 96 -637 98 -633
rect -318 -678 -316 -675
rect -284 -678 -282 -675
rect -249 -677 -247 -674
rect -214 -678 -212 -675
rect -177 -677 -175 -674
rect -140 -676 -138 -673
rect -104 -676 -102 -673
rect -68 -676 -66 -673
rect -34 -675 -32 -672
rect 5 -674 7 -671
rect -318 -794 -316 -778
rect -284 -794 -282 -778
rect -249 -793 -247 -777
rect 174 -716 176 -713
rect 212 -716 214 -713
rect 256 -716 258 -713
rect 294 -716 296 -713
rect 174 -774 176 -756
rect 212 -774 214 -756
rect 256 -774 258 -756
rect 294 -774 296 -756
rect -214 -794 -212 -778
rect -177 -793 -175 -777
rect -140 -792 -138 -776
rect -104 -792 -102 -776
rect -68 -792 -66 -776
rect -34 -791 -32 -775
rect 5 -790 7 -774
rect 174 -798 176 -794
rect 212 -798 214 -794
rect 256 -798 258 -794
rect 294 -798 296 -794
<< metal1 >>
rect 91 -545 95 -542
rect -257 -557 -253 -548
rect -207 -556 -203 -547
rect -157 -556 -153 -547
rect -110 -556 -106 -547
rect 85 -549 86 -545
rect 90 -549 95 -545
rect 91 -555 95 -549
rect -263 -562 -262 -557
rect -258 -562 -239 -557
rect -213 -561 -212 -556
rect -208 -561 -189 -556
rect -163 -561 -162 -556
rect -158 -561 -139 -556
rect -116 -561 -115 -556
rect -111 -561 -92 -556
rect -257 -568 -253 -562
rect -207 -567 -203 -561
rect -157 -567 -153 -561
rect -110 -567 -106 -561
rect 99 -613 103 -595
rect -249 -632 -245 -618
rect -199 -631 -195 -617
rect -149 -631 -145 -617
rect -102 -631 -98 -617
rect 91 -643 95 -633
rect -323 -678 -319 -670
rect -289 -678 -285 -670
rect -254 -677 -250 -669
rect -315 -787 -311 -778
rect -281 -787 -277 -778
rect -246 -786 -242 -777
rect -219 -678 -215 -670
rect -182 -677 -178 -669
rect -145 -676 -141 -668
rect -109 -676 -105 -668
rect -73 -676 -69 -668
rect -39 -675 -35 -667
rect 0 -674 4 -666
rect 169 -706 173 -703
rect 207 -706 211 -703
rect 251 -706 255 -703
rect 289 -706 293 -703
rect 163 -710 164 -706
rect 168 -710 173 -706
rect 201 -710 202 -706
rect 206 -710 211 -706
rect 245 -710 246 -706
rect 250 -710 255 -706
rect 283 -710 284 -706
rect 288 -710 293 -706
rect 169 -716 173 -710
rect 207 -716 211 -710
rect 251 -716 255 -710
rect 289 -716 293 -710
rect 177 -774 181 -756
rect 215 -774 219 -756
rect 259 -774 263 -756
rect 297 -774 301 -756
rect -211 -787 -207 -778
rect -174 -786 -170 -777
rect -137 -785 -133 -776
rect -101 -785 -97 -776
rect -65 -785 -61 -776
rect -31 -784 -27 -775
rect 8 -783 12 -774
rect 169 -804 173 -794
rect 207 -804 211 -794
rect 251 -804 255 -794
rect 289 -804 293 -794
<< pm12contact >>
rect 91 -610 96 -605
rect -258 -641 -252 -635
rect -208 -640 -202 -634
rect -158 -640 -152 -634
rect -111 -640 -105 -634
rect 169 -771 174 -766
rect 207 -771 212 -766
rect 251 -771 256 -766
rect 289 -771 294 -766
rect -323 -794 -318 -789
rect -289 -794 -284 -789
rect -254 -793 -249 -788
rect -219 -794 -214 -789
rect -182 -793 -177 -788
rect -145 -792 -140 -787
rect -109 -792 -104 -787
rect -73 -792 -68 -787
rect -39 -791 -34 -786
rect 0 -790 5 -785
<< metal2 >>
rect 88 -610 91 -605
rect -268 -641 -258 -635
rect -218 -640 -208 -634
rect -168 -640 -158 -634
rect -121 -640 -111 -634
rect 166 -771 169 -766
rect 204 -771 207 -766
rect 248 -771 251 -766
rect 286 -771 289 -766
rect -331 -794 -323 -789
rect -297 -794 -289 -789
rect -262 -793 -254 -788
rect -227 -794 -219 -789
rect -190 -793 -182 -788
rect -153 -792 -145 -787
rect -117 -792 -109 -787
rect -81 -792 -73 -787
rect -47 -791 -39 -786
rect -8 -790 0 -785
<< labels >>
rlabel metal1 -257 -553 -253 -548 5 vdd!
rlabel metal1 -207 -552 -203 -547 5 vdd!
rlabel metal1 -157 -552 -153 -547 5 vdd!
rlabel metal1 -110 -552 -106 -547 5 vdd!
rlabel metal2 -268 -641 -262 -635 2 clock_in
rlabel metal2 -218 -640 -212 -634 1 clock_in
rlabel metal2 -168 -640 -162 -634 1 clock_in
rlabel metal2 -121 -640 -116 -634 1 clock_in
rlabel metal1 -249 -632 -245 -627 1 pdr1
rlabel metal1 -199 -631 -195 -627 1 pdr2
rlabel metal1 -149 -631 -145 -627 1 pdr3
rlabel metal1 -102 -631 -98 -627 1 pdr4
rlabel metal1 -323 -675 -319 -670 1 pdr1
rlabel metal2 -331 -794 -326 -789 2 prop_1
rlabel metal1 -315 -787 -311 -782 1 prop1_car0
rlabel metal1 -289 -675 -285 -670 1 prop1_car0
rlabel metal2 -297 -794 -293 -789 1 carry_0
rlabel metal1 -281 -787 -277 -782 1 clock_car0
rlabel metal1 -254 -673 -250 -669 1 clock_car0
rlabel metal2 -262 -793 -257 -788 1 clock_in
rlabel metal1 -246 -786 -242 -782 1 gnd!
rlabel metal1 -219 -675 -215 -670 1 pdr2
rlabel metal2 -227 -794 -222 -789 1 prop_2
rlabel metal1 -211 -787 -207 -782 1 pdr1
rlabel metal1 -182 -674 -178 -669 1 pdr1
rlabel metal2 -190 -793 -186 -788 1 gen_1
rlabel metal1 -174 -786 -170 -782 1 clock_car0
rlabel metal1 -145 -673 -141 -668 1 pdr3
rlabel metal2 -153 -792 -149 -787 1 prop_3
rlabel metal1 -137 -785 -133 -781 1 pdr2
rlabel metal1 -109 -673 -105 -668 1 pdr2
rlabel metal2 -117 -792 -113 -787 1 gen_2
rlabel metal1 -101 -785 -97 -780 1 clock_car0
rlabel metal1 -73 -672 -69 -668 1 pdr4
rlabel metal2 -81 -792 -77 -787 1 prop_4
rlabel metal1 -65 -785 -61 -781 1 pdr3
rlabel metal1 -39 -672 -35 -667 1 pdr3
rlabel metal2 -47 -791 -43 -786 1 gen_3
rlabel metal1 -31 -784 -27 -780 1 clock_car0
rlabel metal1 0 -671 4 -666 1 pdr4
rlabel metal2 -8 -790 -4 -785 1 gen_4
rlabel metal1 8 -783 12 -778 7 clock_car0
rlabel metal1 169 -707 173 -703 1 vdd!
rlabel metal1 207 -707 211 -703 1 vdd!
rlabel metal1 251 -706 255 -703 1 vdd!
rlabel metal1 289 -706 293 -703 1 vdd!
rlabel metal1 169 -804 173 -800 1 gnd!
rlabel metal1 207 -804 211 -800 1 gnd!
rlabel metal1 251 -804 255 -800 1 gnd!
rlabel metal1 289 -804 293 -800 1 gnd!
rlabel metal2 166 -771 168 -766 1 pdr1
rlabel metal2 204 -771 206 -766 1 pdr2
rlabel metal2 248 -771 250 -766 1 pdr3
rlabel metal2 286 -771 288 -766 1 pdr4
rlabel metal1 178 -771 181 -767 1 c1
rlabel metal1 216 -771 219 -766 1 c2
rlabel metal1 260 -771 263 -766 1 c3
rlabel metal1 298 -771 301 -766 1 c4
rlabel metal1 91 -546 95 -542 1 vdd!
rlabel metal1 91 -643 95 -639 1 gnd!
rlabel metal2 88 -610 91 -605 1 clk_org
rlabel metal1 100 -610 103 -606 1 clock_in
<< end >>
