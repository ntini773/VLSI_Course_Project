magic
tech scmos
timestamp 1731952909
<< nwell >>
rect -57 67 -20 69
rect -57 12 -19 67
rect -13 12 30 64
<< ntransistor >>
rect -43 -38 -41 -18
rect -33 -38 -31 -18
rect 1 -38 3 -18
rect 11 -38 13 -18
<< ptransistor >>
rect -43 18 -41 58
rect -33 18 -31 58
rect 1 18 3 58
rect 11 18 13 58
<< ndiffusion >>
rect -44 -38 -43 -18
rect -41 -38 -33 -18
rect -31 -38 -30 -18
rect 0 -38 1 -18
rect 3 -38 11 -18
rect 13 -38 14 -18
<< pdiffusion >>
rect -44 18 -43 58
rect -41 18 -39 58
rect -35 18 -33 58
rect -31 18 -30 58
rect 0 18 1 58
rect 3 18 5 58
rect 9 18 11 58
rect 13 18 14 58
<< ndcontact >>
rect -48 -38 -44 -18
rect -30 -38 -26 -18
rect -4 -38 0 -18
rect 14 -38 18 -18
<< pdcontact >>
rect -48 18 -44 58
rect -39 18 -35 58
rect -30 18 -26 58
rect -4 18 0 58
rect 5 18 9 58
rect 14 18 18 58
<< psubstratepcontact >>
rect -16 -45 -8 -41
<< nsubstratencontact >>
rect -49 62 -43 66
rect 22 56 27 61
<< polysilicon >>
rect -43 58 -41 61
rect -33 58 -31 61
rect 1 58 3 61
rect 11 58 13 61
rect -43 14 -41 18
rect -42 9 -41 14
rect -43 -18 -41 9
rect -33 -10 -31 18
rect -33 -18 -31 -14
rect 1 -18 3 18
rect 11 -18 13 18
rect -43 -41 -41 -38
rect -33 -41 -31 -38
rect 1 -41 3 -38
rect 11 -41 13 -38
<< polycontact >>
rect -3 1 1 5
rect 7 -7 11 -3
<< metal1 >>
rect -77 74 -58 75
rect -77 70 25 74
rect -49 66 -44 70
rect -49 60 -44 62
rect -48 58 -44 60
rect -30 58 -26 70
rect -103 32 -101 36
rect -81 32 -66 36
rect -70 5 -66 32
rect -4 64 18 67
rect -4 58 0 64
rect 14 58 18 64
rect -39 14 -35 18
rect -4 14 0 18
rect -39 10 0 14
rect 21 61 25 70
rect 21 56 22 61
rect 5 12 9 18
rect 5 8 22 12
rect -70 1 -3 5
rect -66 -7 7 -3
rect -66 -56 -62 -7
rect 18 -11 22 8
rect -16 -15 22 -11
rect -16 -18 -12 -15
rect -105 -60 -102 -56
rect -82 -60 -62 -56
rect -26 -22 -4 -18
rect -48 -41 -44 -38
rect 14 -41 18 -38
rect -48 -45 -16 -41
rect -8 -45 18 -41
rect -48 -77 -44 -45
rect -77 -81 -74 -77
rect -69 -81 -44 -77
<< m2contact >>
rect -109 31 -103 37
rect -111 -61 -105 -55
<< pnm12contact >>
rect -49 9 -42 14
rect -37 -14 -31 -10
<< metal2 >>
rect -108 26 -104 31
rect -108 22 -59 26
rect -63 13 -59 22
rect -63 9 -49 13
rect -110 -10 -54 -8
rect -110 -12 -37 -10
rect -110 -55 -106 -12
rect -58 -14 -37 -12
rect -58 -15 -54 -14
rect -105 -60 -104 -56
<< m123contact >>
rect -103 68 -97 75
rect -88 7 -82 12
rect -102 -24 -97 -17
rect -74 -82 -69 -77
<< metal3 >>
rect -101 -17 -97 68
rect -86 12 -82 14
rect -86 1 -82 7
rect -86 -3 -70 1
rect -74 -77 -70 -3
use inverter  inverter_0
timestamp 1731871317
transform 1 0 -107 0 1 37
box 6 -28 31 40
use inverter  inverter_1
timestamp 1731871317
transform 1 0 -108 0 1 -55
box 6 -28 31 40
<< labels >>
rlabel metal1 -28 72 -28 72 5 vdd
rlabel metal1 20 3 20 3 7 out
rlabel metal1 -16 -43 -16 -43 1 gnd
<< end >>
