magic
tech scmos
timestamp 1732009470
<< nwell >>
rect 3094 -1100 3127 -1053
rect 3146 -1094 3212 -1052
rect 372 -1246 405 -1199
rect 424 -1240 490 -1198
rect 1313 -1347 1337 -1285
rect 1363 -1346 1387 -1284
rect 1413 -1346 1437 -1284
rect 1460 -1346 1484 -1284
rect 102 -1425 138 -1385
rect 144 -1432 168 -1392
rect 1782 -1568 1806 -1516
rect 1820 -1568 1844 -1516
rect 1864 -1568 1888 -1516
rect 1902 -1568 1926 -1516
rect 1948 -1566 1972 -1514
rect 3150 -1521 3183 -1474
rect 3202 -1515 3268 -1473
rect 413 -1622 446 -1575
rect 465 -1616 531 -1574
rect 104 -1775 140 -1735
rect 146 -1782 170 -1742
rect 438 -1931 471 -1884
rect 490 -1925 556 -1883
rect 3170 -1938 3203 -1891
rect 3222 -1932 3288 -1890
rect 112 -2067 148 -2027
rect 154 -2074 178 -2034
rect 434 -2286 467 -2239
rect 486 -2280 552 -2238
rect 3219 -2324 3252 -2277
rect 3271 -2318 3337 -2276
rect 100 -2433 136 -2393
rect 142 -2440 166 -2400
<< ntransistor >>
rect 3110 -1118 3112 -1108
rect 3159 -1121 3161 -1111
rect 3193 -1121 3195 -1111
rect 388 -1264 390 -1254
rect 437 -1267 439 -1257
rect 471 -1267 473 -1257
rect 113 -1468 115 -1448
rect 124 -1468 126 -1448
rect 155 -1450 157 -1440
rect 429 -1640 431 -1630
rect 1260 -1627 1262 -1527
rect 1288 -1627 1290 -1527
rect 1315 -1627 1317 -1527
rect 1354 -1627 1356 -1527
rect 1382 -1627 1384 -1527
rect 1409 -1627 1411 -1527
rect 1449 -1626 1451 -1526
rect 1477 -1626 1479 -1526
rect 1504 -1626 1506 -1526
rect 1540 -1626 1542 -1526
rect 3166 -1539 3168 -1529
rect 3215 -1542 3217 -1532
rect 3249 -1542 3251 -1532
rect 1793 -1600 1795 -1580
rect 1831 -1600 1833 -1580
rect 1875 -1600 1877 -1580
rect 1913 -1600 1915 -1580
rect 1959 -1598 1961 -1578
rect 478 -1643 480 -1633
rect 512 -1643 514 -1633
rect 115 -1818 117 -1798
rect 126 -1818 128 -1798
rect 157 -1800 159 -1790
rect 454 -1949 456 -1939
rect 503 -1952 505 -1942
rect 537 -1952 539 -1942
rect 3186 -1956 3188 -1946
rect 3235 -1959 3237 -1949
rect 3269 -1959 3271 -1949
rect 123 -2110 125 -2090
rect 134 -2110 136 -2090
rect 165 -2092 167 -2082
rect 450 -2304 452 -2294
rect 499 -2307 501 -2297
rect 533 -2307 535 -2297
rect 3235 -2342 3237 -2332
rect 3284 -2345 3286 -2335
rect 3318 -2345 3320 -2335
rect 111 -2476 113 -2456
rect 122 -2476 124 -2456
rect 153 -2458 155 -2448
<< ptransistor >>
rect 3110 -1088 3112 -1068
rect 3159 -1080 3161 -1060
rect 3193 -1080 3195 -1060
rect 388 -1234 390 -1214
rect 437 -1226 439 -1206
rect 471 -1226 473 -1206
rect 1324 -1341 1326 -1291
rect 1374 -1340 1376 -1290
rect 1424 -1340 1426 -1290
rect 1471 -1340 1473 -1290
rect 113 -1419 115 -1399
rect 124 -1419 126 -1399
rect 155 -1426 157 -1406
rect 3166 -1509 3168 -1489
rect 3215 -1501 3217 -1481
rect 3249 -1501 3251 -1481
rect 429 -1610 431 -1590
rect 478 -1602 480 -1582
rect 512 -1602 514 -1582
rect 1793 -1562 1795 -1522
rect 1831 -1562 1833 -1522
rect 1875 -1562 1877 -1522
rect 1913 -1562 1915 -1522
rect 1959 -1560 1961 -1520
rect 115 -1769 117 -1749
rect 126 -1769 128 -1749
rect 157 -1776 159 -1756
rect 454 -1919 456 -1899
rect 503 -1911 505 -1891
rect 537 -1911 539 -1891
rect 3186 -1926 3188 -1906
rect 3235 -1918 3237 -1898
rect 3269 -1918 3271 -1898
rect 123 -2061 125 -2041
rect 134 -2061 136 -2041
rect 165 -2068 167 -2048
rect 450 -2274 452 -2254
rect 499 -2266 501 -2246
rect 533 -2266 535 -2246
rect 3235 -2312 3237 -2292
rect 3284 -2304 3286 -2284
rect 3318 -2304 3320 -2284
rect 111 -2427 113 -2407
rect 122 -2427 124 -2407
rect 153 -2434 155 -2414
<< ndiffusion >>
rect 3109 -1118 3110 -1108
rect 3112 -1118 3113 -1108
rect 3158 -1121 3159 -1111
rect 3161 -1121 3162 -1111
rect 3192 -1121 3193 -1111
rect 3195 -1121 3196 -1111
rect 387 -1264 388 -1254
rect 390 -1264 391 -1254
rect 436 -1267 437 -1257
rect 439 -1267 440 -1257
rect 470 -1267 471 -1257
rect 473 -1267 474 -1257
rect 112 -1468 113 -1448
rect 115 -1468 124 -1448
rect 126 -1468 127 -1448
rect 154 -1450 155 -1440
rect 157 -1450 158 -1440
rect 428 -1640 429 -1630
rect 431 -1640 432 -1630
rect 1259 -1627 1260 -1527
rect 1262 -1627 1263 -1527
rect 1287 -1627 1288 -1527
rect 1290 -1627 1291 -1527
rect 1314 -1627 1315 -1527
rect 1317 -1627 1318 -1527
rect 1353 -1627 1354 -1527
rect 1356 -1627 1357 -1527
rect 1381 -1627 1382 -1527
rect 1384 -1627 1385 -1527
rect 1408 -1627 1409 -1527
rect 1411 -1627 1412 -1527
rect 1448 -1626 1449 -1526
rect 1451 -1626 1452 -1526
rect 1476 -1626 1477 -1526
rect 1479 -1626 1480 -1526
rect 1503 -1626 1504 -1526
rect 1506 -1626 1507 -1526
rect 1539 -1626 1540 -1526
rect 1542 -1626 1543 -1526
rect 3165 -1539 3166 -1529
rect 3168 -1539 3169 -1529
rect 3214 -1542 3215 -1532
rect 3217 -1542 3218 -1532
rect 3248 -1542 3249 -1532
rect 3251 -1542 3252 -1532
rect 1792 -1600 1793 -1580
rect 1795 -1600 1796 -1580
rect 1830 -1600 1831 -1580
rect 1833 -1600 1834 -1580
rect 1874 -1600 1875 -1580
rect 1877 -1600 1878 -1580
rect 1912 -1600 1913 -1580
rect 1915 -1600 1916 -1580
rect 1958 -1598 1959 -1578
rect 1961 -1598 1962 -1578
rect 477 -1643 478 -1633
rect 480 -1643 481 -1633
rect 511 -1643 512 -1633
rect 514 -1643 515 -1633
rect 114 -1818 115 -1798
rect 117 -1818 126 -1798
rect 128 -1818 129 -1798
rect 156 -1800 157 -1790
rect 159 -1800 160 -1790
rect 453 -1949 454 -1939
rect 456 -1949 457 -1939
rect 502 -1952 503 -1942
rect 505 -1952 506 -1942
rect 536 -1952 537 -1942
rect 539 -1952 540 -1942
rect 3185 -1956 3186 -1946
rect 3188 -1956 3189 -1946
rect 3234 -1959 3235 -1949
rect 3237 -1959 3238 -1949
rect 3268 -1959 3269 -1949
rect 3271 -1959 3272 -1949
rect 122 -2110 123 -2090
rect 125 -2110 134 -2090
rect 136 -2110 137 -2090
rect 164 -2092 165 -2082
rect 167 -2092 168 -2082
rect 449 -2304 450 -2294
rect 452 -2304 453 -2294
rect 498 -2307 499 -2297
rect 501 -2307 502 -2297
rect 532 -2307 533 -2297
rect 535 -2307 536 -2297
rect 3234 -2342 3235 -2332
rect 3237 -2342 3238 -2332
rect 3283 -2345 3284 -2335
rect 3286 -2345 3287 -2335
rect 3317 -2345 3318 -2335
rect 3320 -2345 3321 -2335
rect 110 -2476 111 -2456
rect 113 -2476 122 -2456
rect 124 -2476 125 -2456
rect 152 -2458 153 -2448
rect 155 -2458 156 -2448
<< pdiffusion >>
rect 3109 -1088 3110 -1068
rect 3112 -1088 3113 -1068
rect 3158 -1080 3159 -1060
rect 3161 -1080 3162 -1060
rect 3192 -1080 3193 -1060
rect 3195 -1080 3196 -1060
rect 387 -1234 388 -1214
rect 390 -1234 391 -1214
rect 436 -1226 437 -1206
rect 439 -1226 440 -1206
rect 470 -1226 471 -1206
rect 473 -1226 474 -1206
rect 1323 -1341 1324 -1291
rect 1326 -1341 1327 -1291
rect 1373 -1340 1374 -1290
rect 1376 -1340 1377 -1290
rect 1423 -1340 1424 -1290
rect 1426 -1340 1427 -1290
rect 1470 -1340 1471 -1290
rect 1473 -1340 1474 -1290
rect 112 -1419 113 -1399
rect 115 -1419 119 -1399
rect 123 -1419 124 -1399
rect 126 -1419 127 -1399
rect 154 -1426 155 -1406
rect 157 -1426 158 -1406
rect 3165 -1509 3166 -1489
rect 3168 -1509 3169 -1489
rect 3214 -1501 3215 -1481
rect 3217 -1501 3218 -1481
rect 3248 -1501 3249 -1481
rect 3251 -1501 3252 -1481
rect 428 -1610 429 -1590
rect 431 -1610 432 -1590
rect 477 -1602 478 -1582
rect 480 -1602 481 -1582
rect 511 -1602 512 -1582
rect 514 -1602 515 -1582
rect 1792 -1562 1793 -1522
rect 1795 -1562 1796 -1522
rect 1830 -1562 1831 -1522
rect 1833 -1562 1834 -1522
rect 1874 -1562 1875 -1522
rect 1877 -1562 1878 -1522
rect 1912 -1562 1913 -1522
rect 1915 -1562 1916 -1522
rect 1958 -1560 1959 -1520
rect 1961 -1560 1962 -1520
rect 114 -1769 115 -1749
rect 117 -1769 121 -1749
rect 125 -1769 126 -1749
rect 128 -1769 129 -1749
rect 156 -1776 157 -1756
rect 159 -1776 160 -1756
rect 453 -1919 454 -1899
rect 456 -1919 457 -1899
rect 502 -1911 503 -1891
rect 505 -1911 506 -1891
rect 536 -1911 537 -1891
rect 539 -1911 540 -1891
rect 3185 -1926 3186 -1906
rect 3188 -1926 3189 -1906
rect 3234 -1918 3235 -1898
rect 3237 -1918 3238 -1898
rect 3268 -1918 3269 -1898
rect 3271 -1918 3272 -1898
rect 122 -2061 123 -2041
rect 125 -2061 129 -2041
rect 133 -2061 134 -2041
rect 136 -2061 137 -2041
rect 164 -2068 165 -2048
rect 167 -2068 168 -2048
rect 449 -2274 450 -2254
rect 452 -2274 453 -2254
rect 498 -2266 499 -2246
rect 501 -2266 502 -2246
rect 532 -2266 533 -2246
rect 535 -2266 536 -2246
rect 3234 -2312 3235 -2292
rect 3237 -2312 3238 -2292
rect 3283 -2304 3284 -2284
rect 3286 -2304 3287 -2284
rect 3317 -2304 3318 -2284
rect 3320 -2304 3321 -2284
rect 110 -2427 111 -2407
rect 113 -2427 117 -2407
rect 121 -2427 122 -2407
rect 124 -2427 125 -2407
rect 152 -2434 153 -2414
rect 155 -2434 156 -2414
<< ndcontact >>
rect 3105 -1118 3109 -1108
rect 3113 -1118 3117 -1108
rect 3154 -1121 3158 -1111
rect 3162 -1121 3166 -1111
rect 3188 -1121 3192 -1111
rect 3196 -1121 3200 -1111
rect 383 -1264 387 -1254
rect 391 -1264 395 -1254
rect 432 -1267 436 -1257
rect 440 -1267 444 -1257
rect 466 -1267 470 -1257
rect 474 -1267 478 -1257
rect 108 -1468 112 -1448
rect 127 -1468 131 -1448
rect 150 -1450 154 -1440
rect 158 -1450 162 -1440
rect 424 -1640 428 -1630
rect 432 -1640 436 -1630
rect 1255 -1627 1259 -1527
rect 1263 -1627 1267 -1527
rect 1283 -1627 1287 -1527
rect 1291 -1627 1295 -1527
rect 1310 -1627 1314 -1527
rect 1318 -1627 1322 -1527
rect 1349 -1627 1353 -1527
rect 1357 -1627 1361 -1527
rect 1377 -1627 1381 -1527
rect 1385 -1627 1389 -1527
rect 1404 -1627 1408 -1527
rect 1412 -1627 1416 -1527
rect 1444 -1626 1448 -1526
rect 1452 -1626 1456 -1526
rect 1472 -1626 1476 -1526
rect 1480 -1626 1484 -1526
rect 1499 -1626 1503 -1526
rect 1507 -1626 1511 -1526
rect 1535 -1626 1539 -1526
rect 1543 -1626 1547 -1526
rect 3161 -1539 3165 -1529
rect 3169 -1539 3173 -1529
rect 3210 -1542 3214 -1532
rect 3218 -1542 3222 -1532
rect 3244 -1542 3248 -1532
rect 3252 -1542 3256 -1532
rect 1788 -1600 1792 -1580
rect 1796 -1600 1800 -1580
rect 1826 -1600 1830 -1580
rect 1834 -1600 1838 -1580
rect 1870 -1600 1874 -1580
rect 1878 -1600 1882 -1580
rect 1908 -1600 1912 -1580
rect 1916 -1600 1920 -1580
rect 1954 -1598 1958 -1578
rect 1962 -1598 1966 -1578
rect 473 -1643 477 -1633
rect 481 -1643 485 -1633
rect 507 -1643 511 -1633
rect 515 -1643 519 -1633
rect 110 -1818 114 -1798
rect 129 -1818 133 -1798
rect 152 -1800 156 -1790
rect 160 -1800 164 -1790
rect 449 -1949 453 -1939
rect 457 -1949 461 -1939
rect 498 -1952 502 -1942
rect 506 -1952 510 -1942
rect 532 -1952 536 -1942
rect 540 -1952 544 -1942
rect 3181 -1956 3185 -1946
rect 3189 -1956 3193 -1946
rect 3230 -1959 3234 -1949
rect 3238 -1959 3242 -1949
rect 3264 -1959 3268 -1949
rect 3272 -1959 3276 -1949
rect 118 -2110 122 -2090
rect 137 -2110 141 -2090
rect 160 -2092 164 -2082
rect 168 -2092 172 -2082
rect 445 -2304 449 -2294
rect 453 -2304 457 -2294
rect 494 -2307 498 -2297
rect 502 -2307 506 -2297
rect 528 -2307 532 -2297
rect 536 -2307 540 -2297
rect 3230 -2342 3234 -2332
rect 3238 -2342 3242 -2332
rect 3279 -2345 3283 -2335
rect 3287 -2345 3291 -2335
rect 3313 -2345 3317 -2335
rect 3321 -2345 3325 -2335
rect 106 -2476 110 -2456
rect 125 -2476 129 -2456
rect 148 -2458 152 -2448
rect 156 -2458 160 -2448
<< pdcontact >>
rect 3105 -1088 3109 -1068
rect 3113 -1088 3117 -1068
rect 3154 -1080 3158 -1060
rect 3162 -1080 3166 -1060
rect 3188 -1080 3192 -1060
rect 3196 -1080 3200 -1060
rect 383 -1234 387 -1214
rect 391 -1234 395 -1214
rect 432 -1226 436 -1206
rect 440 -1226 444 -1206
rect 466 -1226 470 -1206
rect 474 -1226 478 -1206
rect 1319 -1341 1323 -1291
rect 1327 -1341 1331 -1291
rect 1369 -1340 1373 -1290
rect 1377 -1340 1381 -1290
rect 1419 -1340 1423 -1290
rect 1427 -1340 1431 -1290
rect 1466 -1340 1470 -1290
rect 1474 -1340 1478 -1290
rect 108 -1419 112 -1399
rect 119 -1419 123 -1399
rect 127 -1419 131 -1399
rect 150 -1426 154 -1406
rect 158 -1426 162 -1406
rect 3161 -1509 3165 -1489
rect 3169 -1509 3173 -1489
rect 3210 -1501 3214 -1481
rect 3218 -1501 3222 -1481
rect 3244 -1501 3248 -1481
rect 3252 -1501 3256 -1481
rect 424 -1610 428 -1590
rect 432 -1610 436 -1590
rect 473 -1602 477 -1582
rect 481 -1602 485 -1582
rect 507 -1602 511 -1582
rect 515 -1602 519 -1582
rect 1788 -1562 1792 -1522
rect 1796 -1562 1800 -1522
rect 1826 -1562 1830 -1522
rect 1834 -1562 1838 -1522
rect 1870 -1562 1874 -1522
rect 1878 -1562 1882 -1522
rect 1908 -1562 1912 -1522
rect 1916 -1562 1920 -1522
rect 1954 -1560 1958 -1520
rect 1962 -1560 1966 -1520
rect 110 -1769 114 -1749
rect 121 -1769 125 -1749
rect 129 -1769 133 -1749
rect 152 -1776 156 -1756
rect 160 -1776 164 -1756
rect 449 -1919 453 -1899
rect 457 -1919 461 -1899
rect 498 -1911 502 -1891
rect 506 -1911 510 -1891
rect 532 -1911 536 -1891
rect 540 -1911 544 -1891
rect 3181 -1926 3185 -1906
rect 3189 -1926 3193 -1906
rect 3230 -1918 3234 -1898
rect 3238 -1918 3242 -1898
rect 3264 -1918 3268 -1898
rect 3272 -1918 3276 -1898
rect 118 -2061 122 -2041
rect 129 -2061 133 -2041
rect 137 -2061 141 -2041
rect 160 -2068 164 -2048
rect 168 -2068 172 -2048
rect 445 -2274 449 -2254
rect 453 -2274 457 -2254
rect 494 -2266 498 -2246
rect 502 -2266 506 -2246
rect 528 -2266 532 -2246
rect 536 -2266 540 -2246
rect 3230 -2312 3234 -2292
rect 3238 -2312 3242 -2292
rect 3279 -2304 3283 -2284
rect 3287 -2304 3291 -2284
rect 3313 -2304 3317 -2284
rect 3321 -2304 3325 -2284
rect 106 -2427 110 -2407
rect 117 -2427 121 -2407
rect 125 -2427 129 -2407
rect 148 -2434 152 -2414
rect 156 -2434 160 -2414
<< psubstratepcontact >>
rect 164 -1459 169 -1455
rect 166 -1809 171 -1805
rect 174 -2101 179 -2097
rect 162 -2467 167 -2463
<< nsubstratencontact >>
rect 1314 -1285 1318 -1280
rect 1364 -1284 1368 -1279
rect 1414 -1284 1418 -1279
rect 1461 -1284 1465 -1279
rect 108 -1394 112 -1388
rect 160 -1399 164 -1395
rect 1783 -1516 1787 -1512
rect 1821 -1516 1825 -1512
rect 1865 -1516 1869 -1512
rect 1903 -1516 1907 -1512
rect 1949 -1514 1953 -1510
rect 110 -1744 114 -1738
rect 162 -1749 166 -1745
rect 118 -2036 122 -2030
rect 170 -2041 174 -2037
rect 106 -2402 110 -2396
rect 158 -2407 162 -2403
<< polysilicon >>
rect 3110 -1068 3112 -1059
rect 3159 -1060 3161 -1053
rect 3193 -1060 3195 -1056
rect 3110 -1108 3112 -1088
rect 3159 -1095 3161 -1080
rect 3159 -1111 3161 -1108
rect 3193 -1111 3195 -1080
rect 3110 -1121 3112 -1118
rect 3159 -1140 3161 -1121
rect 3193 -1124 3195 -1121
rect 388 -1214 390 -1205
rect 437 -1206 439 -1199
rect 471 -1206 473 -1202
rect 388 -1254 390 -1234
rect 437 -1241 439 -1226
rect 437 -1257 439 -1254
rect 471 -1257 473 -1226
rect 388 -1267 390 -1264
rect 437 -1286 439 -1267
rect 471 -1270 473 -1267
rect 1324 -1291 1326 -1288
rect 1374 -1290 1376 -1287
rect 1424 -1290 1426 -1287
rect 1471 -1290 1473 -1287
rect 1324 -1364 1326 -1341
rect 1374 -1363 1376 -1340
rect 1424 -1363 1426 -1340
rect 1471 -1363 1473 -1340
rect 113 -1399 115 -1396
rect 124 -1399 126 -1396
rect 155 -1406 157 -1402
rect 113 -1448 115 -1419
rect 124 -1448 126 -1419
rect 155 -1440 157 -1426
rect 155 -1453 157 -1450
rect 113 -1471 115 -1468
rect 124 -1471 126 -1468
rect 3166 -1489 3168 -1480
rect 3215 -1481 3217 -1474
rect 3249 -1481 3251 -1477
rect 1793 -1522 1795 -1519
rect 1831 -1522 1833 -1519
rect 1875 -1522 1877 -1519
rect 1913 -1522 1915 -1519
rect 1959 -1520 1961 -1517
rect 1260 -1527 1262 -1524
rect 1288 -1527 1290 -1524
rect 1315 -1527 1317 -1524
rect 1354 -1527 1356 -1524
rect 1382 -1527 1384 -1524
rect 1409 -1527 1411 -1524
rect 1449 -1526 1451 -1523
rect 1477 -1526 1479 -1523
rect 1504 -1526 1506 -1523
rect 1540 -1526 1542 -1523
rect 429 -1590 431 -1581
rect 478 -1582 480 -1575
rect 512 -1582 514 -1578
rect 429 -1630 431 -1610
rect 478 -1617 480 -1602
rect 478 -1633 480 -1630
rect 512 -1633 514 -1602
rect 3166 -1529 3168 -1509
rect 3215 -1516 3217 -1501
rect 3215 -1532 3217 -1529
rect 3249 -1532 3251 -1501
rect 3166 -1542 3168 -1539
rect 1793 -1580 1795 -1562
rect 1831 -1580 1833 -1562
rect 1875 -1580 1877 -1562
rect 1913 -1580 1915 -1562
rect 1959 -1578 1961 -1560
rect 3215 -1561 3217 -1542
rect 3249 -1545 3251 -1542
rect 1793 -1604 1795 -1600
rect 1831 -1604 1833 -1600
rect 1875 -1604 1877 -1600
rect 1913 -1604 1915 -1600
rect 1959 -1602 1961 -1598
rect 429 -1643 431 -1640
rect 1260 -1639 1262 -1627
rect 1288 -1639 1290 -1627
rect 1315 -1639 1317 -1627
rect 1354 -1639 1356 -1627
rect 1382 -1639 1384 -1627
rect 1409 -1639 1411 -1627
rect 1449 -1638 1451 -1626
rect 1477 -1638 1479 -1626
rect 1504 -1638 1506 -1626
rect 1540 -1638 1542 -1626
rect 478 -1662 480 -1643
rect 512 -1646 514 -1643
rect 115 -1749 117 -1746
rect 126 -1749 128 -1746
rect 157 -1756 159 -1752
rect 115 -1798 117 -1769
rect 126 -1798 128 -1769
rect 157 -1790 159 -1776
rect 157 -1803 159 -1800
rect 115 -1821 117 -1818
rect 126 -1821 128 -1818
rect 454 -1899 456 -1890
rect 503 -1891 505 -1884
rect 537 -1891 539 -1887
rect 3186 -1906 3188 -1897
rect 3235 -1898 3237 -1891
rect 3269 -1898 3271 -1894
rect 454 -1939 456 -1919
rect 503 -1926 505 -1911
rect 503 -1942 505 -1939
rect 537 -1942 539 -1911
rect 454 -1952 456 -1949
rect 3186 -1946 3188 -1926
rect 3235 -1933 3237 -1918
rect 503 -1971 505 -1952
rect 537 -1955 539 -1952
rect 3235 -1949 3237 -1946
rect 3269 -1949 3271 -1918
rect 3186 -1959 3188 -1956
rect 3235 -1978 3237 -1959
rect 3269 -1962 3271 -1959
rect 123 -2041 125 -2038
rect 134 -2041 136 -2038
rect 165 -2048 167 -2044
rect 123 -2090 125 -2061
rect 134 -2090 136 -2061
rect 165 -2082 167 -2068
rect 165 -2095 167 -2092
rect 123 -2113 125 -2110
rect 134 -2113 136 -2110
rect 450 -2254 452 -2245
rect 499 -2246 501 -2239
rect 533 -2246 535 -2242
rect 450 -2294 452 -2274
rect 499 -2281 501 -2266
rect 499 -2297 501 -2294
rect 533 -2297 535 -2266
rect 3235 -2292 3237 -2283
rect 3284 -2284 3286 -2277
rect 3318 -2284 3320 -2280
rect 450 -2307 452 -2304
rect 499 -2326 501 -2307
rect 533 -2310 535 -2307
rect 3235 -2332 3237 -2312
rect 3284 -2319 3286 -2304
rect 3284 -2335 3286 -2332
rect 3318 -2335 3320 -2304
rect 3235 -2345 3237 -2342
rect 3284 -2364 3286 -2345
rect 3318 -2348 3320 -2345
rect 111 -2407 113 -2404
rect 122 -2407 124 -2404
rect 153 -2414 155 -2410
rect 111 -2456 113 -2427
rect 122 -2456 124 -2427
rect 153 -2448 155 -2434
rect 153 -2461 155 -2458
rect 111 -2479 113 -2476
rect 122 -2479 124 -2476
<< polycontact >>
rect 3161 -1057 3165 -1053
rect 3106 -1105 3110 -1101
rect 3189 -1104 3193 -1100
rect 3161 -1140 3166 -1135
rect 439 -1203 443 -1199
rect 384 -1251 388 -1247
rect 467 -1250 471 -1246
rect 439 -1286 444 -1281
rect 109 -1445 113 -1441
rect 120 -1438 124 -1434
rect 151 -1437 155 -1433
rect 3217 -1478 3221 -1474
rect 480 -1579 484 -1575
rect 425 -1627 429 -1623
rect 508 -1626 512 -1622
rect 3162 -1526 3166 -1522
rect 3245 -1525 3249 -1521
rect 3217 -1561 3222 -1556
rect 480 -1662 485 -1657
rect 111 -1795 115 -1791
rect 122 -1788 126 -1784
rect 153 -1787 157 -1783
rect 505 -1888 509 -1884
rect 3237 -1895 3241 -1891
rect 450 -1936 454 -1932
rect 533 -1935 537 -1931
rect 3182 -1943 3186 -1939
rect 3265 -1942 3269 -1938
rect 505 -1971 510 -1966
rect 3237 -1978 3242 -1973
rect 119 -2087 123 -2083
rect 130 -2080 134 -2076
rect 161 -2079 165 -2075
rect 501 -2243 505 -2239
rect 446 -2291 450 -2287
rect 529 -2290 533 -2286
rect 3286 -2281 3290 -2277
rect 501 -2326 506 -2321
rect 3231 -2329 3235 -2325
rect 3314 -2328 3318 -2324
rect 3286 -2364 3291 -2359
rect 107 -2453 111 -2449
rect 118 -2446 122 -2442
rect 149 -2445 153 -2441
<< metal1 >>
rect 3137 -1030 3144 -1021
rect 3171 -1039 3178 -1023
rect 3079 -1043 3178 -1039
rect 3079 -1101 3088 -1043
rect 3094 -1053 3137 -1046
rect 3171 -1053 3178 -1043
rect 3105 -1068 3109 -1053
rect 3165 -1057 3192 -1053
rect 3188 -1060 3192 -1057
rect 3079 -1105 3106 -1101
rect 3113 -1102 3117 -1088
rect 3154 -1099 3158 -1080
rect 3113 -1106 3140 -1102
rect 3113 -1108 3117 -1106
rect 3105 -1123 3109 -1118
rect 3094 -1130 3130 -1123
rect 3135 -1144 3140 -1106
rect 3154 -1111 3158 -1105
rect 3154 -1127 3158 -1121
rect 3162 -1111 3166 -1080
rect 3196 -1099 3200 -1080
rect 3182 -1104 3189 -1100
rect 3196 -1105 3220 -1099
rect 3196 -1111 3200 -1105
rect 3183 -1117 3188 -1111
rect 3162 -1128 3166 -1121
rect 3196 -1128 3200 -1121
rect 3162 -1132 3200 -1128
rect 3166 -1140 3170 -1135
rect 3135 -1152 3176 -1144
rect 415 -1176 422 -1167
rect 449 -1185 456 -1169
rect 3153 -1176 3158 -1164
rect 357 -1189 456 -1185
rect 357 -1247 366 -1189
rect 372 -1199 415 -1192
rect 449 -1199 456 -1189
rect 383 -1214 387 -1199
rect 443 -1203 470 -1199
rect 466 -1206 470 -1203
rect 357 -1251 384 -1247
rect 391 -1248 395 -1234
rect 432 -1245 436 -1226
rect 391 -1252 418 -1248
rect 391 -1254 395 -1252
rect 383 -1269 387 -1264
rect 372 -1276 408 -1269
rect 413 -1290 418 -1252
rect 432 -1257 436 -1251
rect 432 -1273 436 -1267
rect 440 -1257 444 -1226
rect 474 -1245 478 -1226
rect 460 -1250 467 -1246
rect 474 -1251 498 -1245
rect 474 -1257 478 -1251
rect 461 -1263 466 -1257
rect 440 -1274 444 -1267
rect 474 -1274 478 -1267
rect 440 -1278 478 -1274
rect 1319 -1280 1323 -1271
rect 1369 -1279 1373 -1270
rect 1419 -1279 1423 -1270
rect 1466 -1279 1470 -1270
rect 444 -1286 448 -1281
rect 1313 -1285 1314 -1280
rect 1318 -1285 1337 -1280
rect 1363 -1284 1364 -1279
rect 1368 -1284 1387 -1279
rect 1413 -1284 1414 -1279
rect 1418 -1284 1437 -1279
rect 1460 -1284 1461 -1279
rect 1465 -1284 1484 -1279
rect 413 -1298 454 -1290
rect 1319 -1291 1323 -1285
rect 1369 -1290 1373 -1284
rect 1419 -1290 1423 -1284
rect 1466 -1290 1470 -1284
rect 431 -1322 436 -1310
rect 1327 -1355 1331 -1341
rect 1377 -1354 1381 -1340
rect 1427 -1354 1431 -1340
rect 1474 -1354 1478 -1340
rect 108 -1388 131 -1384
rect 112 -1390 131 -1388
rect 108 -1399 112 -1394
rect 127 -1399 131 -1390
rect 144 -1395 168 -1394
rect 144 -1399 160 -1395
rect 164 -1399 168 -1395
rect 144 -1401 168 -1399
rect 150 -1406 154 -1401
rect 119 -1427 123 -1419
rect 119 -1431 131 -1427
rect 127 -1433 131 -1431
rect 158 -1433 162 -1426
rect 102 -1438 120 -1434
rect 127 -1437 151 -1433
rect 158 -1437 168 -1433
rect 102 -1445 109 -1441
rect 127 -1448 131 -1437
rect 158 -1440 162 -1437
rect 150 -1454 154 -1450
rect 3193 -1451 3200 -1442
rect 144 -1455 169 -1454
rect 144 -1459 164 -1455
rect 144 -1460 169 -1459
rect 3227 -1460 3234 -1444
rect 3135 -1464 3234 -1460
rect 108 -1472 112 -1468
rect 108 -1476 124 -1472
rect 1788 -1509 1808 -1505
rect 1819 -1509 1850 -1505
rect 1862 -1509 1890 -1505
rect 1900 -1509 1921 -1505
rect 1937 -1507 1967 -1503
rect 1788 -1512 1792 -1509
rect 1826 -1512 1830 -1509
rect 1870 -1512 1874 -1509
rect 1908 -1512 1912 -1509
rect 1954 -1510 1958 -1507
rect 1782 -1516 1783 -1512
rect 1787 -1516 1792 -1512
rect 1820 -1516 1821 -1512
rect 1825 -1516 1830 -1512
rect 1864 -1516 1865 -1512
rect 1869 -1516 1874 -1512
rect 1902 -1516 1903 -1512
rect 1907 -1516 1912 -1512
rect 1948 -1514 1949 -1510
rect 1953 -1514 1958 -1510
rect 1255 -1527 1259 -1519
rect 1283 -1527 1287 -1519
rect 1310 -1527 1314 -1519
rect 1349 -1527 1353 -1519
rect 1377 -1527 1381 -1519
rect 1404 -1527 1408 -1519
rect 1444 -1526 1448 -1518
rect 1472 -1526 1476 -1518
rect 1499 -1526 1503 -1518
rect 1535 -1526 1539 -1518
rect 1788 -1522 1792 -1516
rect 1826 -1522 1830 -1516
rect 1870 -1522 1874 -1516
rect 1908 -1522 1912 -1516
rect 1954 -1520 1958 -1514
rect 456 -1552 463 -1543
rect 490 -1561 497 -1545
rect 398 -1565 497 -1561
rect 398 -1623 407 -1565
rect 413 -1575 456 -1568
rect 490 -1575 497 -1565
rect 424 -1590 428 -1575
rect 484 -1579 511 -1575
rect 507 -1582 511 -1579
rect 398 -1627 425 -1623
rect 432 -1624 436 -1610
rect 473 -1621 477 -1602
rect 432 -1628 459 -1624
rect 432 -1630 436 -1628
rect 424 -1645 428 -1640
rect 413 -1652 449 -1645
rect 454 -1666 459 -1628
rect 473 -1633 477 -1627
rect 473 -1649 477 -1643
rect 481 -1633 485 -1602
rect 515 -1621 519 -1602
rect 501 -1626 508 -1622
rect 515 -1627 539 -1621
rect 3135 -1522 3144 -1464
rect 3150 -1474 3193 -1467
rect 3227 -1474 3234 -1464
rect 3161 -1489 3165 -1474
rect 3221 -1478 3248 -1474
rect 3244 -1481 3248 -1478
rect 3135 -1526 3162 -1522
rect 3169 -1523 3173 -1509
rect 3210 -1520 3214 -1501
rect 3169 -1527 3196 -1523
rect 3169 -1529 3173 -1527
rect 3161 -1544 3165 -1539
rect 3150 -1551 3186 -1544
rect 1796 -1580 1800 -1562
rect 1834 -1580 1838 -1562
rect 1878 -1580 1882 -1562
rect 1916 -1580 1920 -1562
rect 1962 -1578 1966 -1560
rect 3191 -1565 3196 -1527
rect 3210 -1532 3214 -1526
rect 3210 -1548 3214 -1542
rect 3218 -1532 3222 -1501
rect 3252 -1520 3256 -1501
rect 3238 -1525 3245 -1521
rect 3252 -1526 3276 -1520
rect 3252 -1532 3256 -1526
rect 3239 -1538 3244 -1532
rect 3218 -1549 3222 -1542
rect 3252 -1549 3256 -1542
rect 3218 -1553 3256 -1549
rect 3222 -1561 3226 -1556
rect 3191 -1573 3232 -1565
rect 3209 -1597 3214 -1585
rect 1788 -1609 1792 -1600
rect 1826 -1609 1830 -1600
rect 1870 -1609 1874 -1600
rect 1908 -1609 1912 -1600
rect 1954 -1607 1958 -1598
rect 1788 -1613 1808 -1609
rect 1819 -1613 1850 -1609
rect 1862 -1613 1890 -1609
rect 1900 -1613 1917 -1609
rect 1937 -1611 1963 -1607
rect 515 -1633 519 -1627
rect 1263 -1633 1267 -1627
rect 1291 -1633 1295 -1627
rect 1318 -1633 1322 -1627
rect 1357 -1633 1361 -1627
rect 1385 -1633 1389 -1627
rect 1412 -1633 1416 -1627
rect 1452 -1632 1456 -1626
rect 1480 -1632 1484 -1626
rect 1507 -1632 1511 -1626
rect 1543 -1632 1547 -1626
rect 502 -1639 507 -1633
rect 481 -1650 485 -1643
rect 515 -1650 519 -1643
rect 481 -1654 519 -1650
rect 485 -1662 489 -1657
rect 454 -1674 495 -1666
rect 472 -1698 477 -1686
rect 110 -1738 133 -1734
rect 114 -1740 133 -1738
rect 110 -1749 114 -1744
rect 129 -1749 133 -1740
rect 146 -1745 170 -1744
rect 146 -1749 162 -1745
rect 166 -1749 170 -1745
rect 146 -1751 170 -1749
rect 152 -1756 156 -1751
rect 121 -1777 125 -1769
rect 121 -1781 133 -1777
rect 129 -1783 133 -1781
rect 160 -1783 164 -1776
rect 104 -1788 122 -1784
rect 129 -1787 153 -1783
rect 160 -1787 170 -1783
rect 104 -1795 111 -1791
rect 129 -1798 133 -1787
rect 160 -1790 164 -1787
rect 152 -1804 156 -1800
rect 146 -1805 171 -1804
rect 146 -1809 166 -1805
rect 146 -1810 171 -1809
rect 110 -1822 114 -1818
rect 110 -1826 126 -1822
rect 481 -1861 488 -1852
rect 515 -1870 522 -1854
rect 423 -1874 522 -1870
rect 3213 -1868 3220 -1859
rect 423 -1932 432 -1874
rect 438 -1884 481 -1877
rect 515 -1884 522 -1874
rect 3247 -1877 3254 -1861
rect 3155 -1881 3254 -1877
rect 449 -1899 453 -1884
rect 509 -1888 536 -1884
rect 532 -1891 536 -1888
rect 423 -1936 450 -1932
rect 457 -1933 461 -1919
rect 498 -1930 502 -1911
rect 457 -1937 484 -1933
rect 457 -1939 461 -1937
rect 449 -1954 453 -1949
rect 438 -1961 474 -1954
rect 479 -1975 484 -1937
rect 498 -1942 502 -1936
rect 498 -1958 502 -1952
rect 506 -1942 510 -1911
rect 540 -1930 544 -1911
rect 526 -1935 533 -1931
rect 540 -1936 564 -1930
rect 540 -1942 544 -1936
rect 527 -1948 532 -1942
rect 3155 -1939 3164 -1881
rect 3170 -1891 3213 -1884
rect 3247 -1891 3254 -1881
rect 3181 -1906 3185 -1891
rect 3241 -1895 3268 -1891
rect 3264 -1898 3268 -1895
rect 3155 -1943 3182 -1939
rect 3189 -1940 3193 -1926
rect 3230 -1937 3234 -1918
rect 3189 -1944 3216 -1940
rect 3189 -1946 3193 -1944
rect 506 -1959 510 -1952
rect 540 -1959 544 -1952
rect 506 -1963 544 -1959
rect 3181 -1961 3185 -1956
rect 510 -1971 514 -1966
rect 3170 -1968 3206 -1961
rect 479 -1983 520 -1975
rect 3211 -1982 3216 -1944
rect 3230 -1949 3234 -1943
rect 3230 -1965 3234 -1959
rect 3238 -1949 3242 -1918
rect 3272 -1937 3276 -1918
rect 3258 -1942 3265 -1938
rect 3272 -1943 3296 -1937
rect 3272 -1949 3276 -1943
rect 3259 -1955 3264 -1949
rect 3238 -1966 3242 -1959
rect 3272 -1966 3276 -1959
rect 3238 -1970 3276 -1966
rect 3242 -1978 3246 -1973
rect 3211 -1990 3252 -1982
rect 497 -2007 502 -1995
rect 3229 -2014 3234 -2002
rect 118 -2030 141 -2026
rect 122 -2032 141 -2030
rect 118 -2041 122 -2036
rect 137 -2041 141 -2032
rect 154 -2037 178 -2036
rect 154 -2041 170 -2037
rect 174 -2041 178 -2037
rect 154 -2043 178 -2041
rect 160 -2048 164 -2043
rect 129 -2069 133 -2061
rect 129 -2073 141 -2069
rect 137 -2075 141 -2073
rect 168 -2075 172 -2068
rect 112 -2080 130 -2076
rect 137 -2079 161 -2075
rect 168 -2079 178 -2075
rect 112 -2087 119 -2083
rect 137 -2090 141 -2079
rect 168 -2082 172 -2079
rect 160 -2096 164 -2092
rect 154 -2097 179 -2096
rect 154 -2101 174 -2097
rect 154 -2102 179 -2101
rect 118 -2114 122 -2110
rect 118 -2118 134 -2114
rect 477 -2216 484 -2207
rect 511 -2225 518 -2209
rect 419 -2229 518 -2225
rect 419 -2287 428 -2229
rect 434 -2239 477 -2232
rect 511 -2239 518 -2229
rect 445 -2254 449 -2239
rect 505 -2243 532 -2239
rect 528 -2246 532 -2243
rect 419 -2291 446 -2287
rect 453 -2288 457 -2274
rect 494 -2285 498 -2266
rect 3262 -2254 3269 -2245
rect 3296 -2263 3303 -2247
rect 453 -2292 480 -2288
rect 453 -2294 457 -2292
rect 445 -2309 449 -2304
rect 434 -2316 470 -2309
rect 475 -2330 480 -2292
rect 494 -2297 498 -2291
rect 494 -2313 498 -2307
rect 502 -2297 506 -2266
rect 536 -2285 540 -2266
rect 3204 -2267 3303 -2263
rect 522 -2290 529 -2286
rect 536 -2291 560 -2285
rect 536 -2297 540 -2291
rect 523 -2303 528 -2297
rect 502 -2314 506 -2307
rect 536 -2314 540 -2307
rect 502 -2318 540 -2314
rect 506 -2326 510 -2321
rect 3204 -2325 3213 -2267
rect 3219 -2277 3262 -2270
rect 3296 -2277 3303 -2267
rect 3230 -2292 3234 -2277
rect 3290 -2281 3317 -2277
rect 3313 -2284 3317 -2281
rect 3204 -2329 3231 -2325
rect 3238 -2326 3242 -2312
rect 3279 -2323 3283 -2304
rect 3238 -2330 3265 -2326
rect 475 -2338 516 -2330
rect 3238 -2332 3242 -2330
rect 3230 -2347 3234 -2342
rect 493 -2362 498 -2350
rect 3219 -2354 3255 -2347
rect 3260 -2368 3265 -2330
rect 3279 -2335 3283 -2329
rect 3279 -2351 3283 -2345
rect 3287 -2335 3291 -2304
rect 3321 -2323 3325 -2304
rect 3307 -2328 3314 -2324
rect 3321 -2329 3345 -2323
rect 3321 -2335 3325 -2329
rect 3308 -2341 3313 -2335
rect 3287 -2352 3291 -2345
rect 3321 -2352 3325 -2345
rect 3287 -2356 3325 -2352
rect 3291 -2364 3295 -2359
rect 3260 -2376 3301 -2368
rect 106 -2396 129 -2392
rect 110 -2398 129 -2396
rect 106 -2407 110 -2402
rect 125 -2407 129 -2398
rect 3278 -2400 3283 -2388
rect 142 -2403 166 -2402
rect 142 -2407 158 -2403
rect 162 -2407 166 -2403
rect 142 -2409 166 -2407
rect 148 -2414 152 -2409
rect 117 -2435 121 -2427
rect 117 -2439 129 -2435
rect 125 -2441 129 -2439
rect 156 -2441 160 -2434
rect 100 -2446 118 -2442
rect 125 -2445 149 -2441
rect 156 -2445 166 -2441
rect 100 -2453 107 -2449
rect 125 -2456 129 -2445
rect 156 -2448 160 -2445
rect 148 -2462 152 -2458
rect 142 -2463 167 -2462
rect 142 -2467 162 -2463
rect 142 -2468 167 -2467
rect 106 -2480 110 -2476
rect 106 -2484 122 -2480
<< m2contact >>
rect 3137 -1036 3144 -1030
rect 3137 -1053 3144 -1046
rect 3153 -1105 3159 -1099
rect 3153 -1132 3158 -1127
rect 3177 -1105 3182 -1099
rect 3176 -1117 3183 -1111
rect 3170 -1140 3175 -1135
rect 3176 -1152 3183 -1144
rect 3153 -1164 3158 -1158
rect 415 -1182 422 -1176
rect 415 -1199 422 -1192
rect 431 -1251 437 -1245
rect 431 -1278 436 -1273
rect 455 -1251 460 -1245
rect 454 -1263 461 -1257
rect 448 -1286 453 -1281
rect 454 -1298 461 -1290
rect 431 -1310 436 -1304
rect 3193 -1457 3200 -1451
rect 456 -1558 463 -1552
rect 456 -1575 463 -1568
rect 472 -1627 478 -1621
rect 472 -1654 477 -1649
rect 496 -1627 501 -1621
rect 3193 -1474 3200 -1467
rect 3209 -1526 3215 -1520
rect 3209 -1553 3214 -1548
rect 3233 -1526 3238 -1520
rect 3232 -1538 3239 -1532
rect 3226 -1561 3231 -1556
rect 3232 -1573 3239 -1565
rect 3209 -1585 3214 -1579
rect 495 -1639 502 -1633
rect 489 -1662 494 -1657
rect 495 -1674 502 -1666
rect 472 -1686 477 -1680
rect 481 -1867 488 -1861
rect 3213 -1874 3220 -1868
rect 481 -1884 488 -1877
rect 497 -1936 503 -1930
rect 497 -1963 502 -1958
rect 521 -1936 526 -1930
rect 520 -1948 527 -1942
rect 3213 -1891 3220 -1884
rect 3229 -1943 3235 -1937
rect 514 -1971 519 -1966
rect 520 -1983 527 -1975
rect 3229 -1970 3234 -1965
rect 3253 -1943 3258 -1937
rect 3252 -1955 3259 -1949
rect 3246 -1978 3251 -1973
rect 497 -1995 502 -1989
rect 3252 -1990 3259 -1982
rect 3229 -2002 3234 -1996
rect 477 -2222 484 -2216
rect 477 -2239 484 -2232
rect 3262 -2260 3269 -2254
rect 493 -2291 499 -2285
rect 493 -2318 498 -2313
rect 517 -2291 522 -2285
rect 516 -2303 523 -2297
rect 510 -2326 515 -2321
rect 3262 -2277 3269 -2270
rect 3278 -2329 3284 -2323
rect 516 -2338 523 -2330
rect 493 -2350 498 -2344
rect 3278 -2356 3283 -2351
rect 3302 -2329 3307 -2323
rect 3301 -2341 3308 -2335
rect 3295 -2364 3300 -2359
rect 3301 -2376 3308 -2368
rect 3278 -2388 3283 -2382
<< pm12contact >>
rect 1318 -1364 1324 -1358
rect 1368 -1363 1374 -1357
rect 1418 -1363 1424 -1357
rect 1465 -1363 1471 -1357
rect 1788 -1577 1793 -1572
rect 1826 -1577 1831 -1572
rect 1870 -1577 1875 -1572
rect 1908 -1577 1913 -1572
rect 1954 -1575 1959 -1570
rect 1255 -1639 1260 -1634
rect 1283 -1639 1288 -1634
rect 1310 -1639 1315 -1634
rect 1349 -1639 1354 -1634
rect 1377 -1639 1382 -1634
rect 1404 -1639 1409 -1634
rect 1444 -1638 1449 -1633
rect 1472 -1638 1477 -1633
rect 1499 -1638 1504 -1633
rect 1535 -1638 1540 -1633
<< metal2 >>
rect 3137 -1046 3144 -1036
rect 3159 -1104 3177 -1100
rect 3153 -1158 3158 -1132
rect 3176 -1135 3183 -1117
rect 3175 -1140 3183 -1135
rect 3176 -1144 3183 -1140
rect 415 -1192 422 -1182
rect 437 -1250 455 -1246
rect 431 -1304 436 -1278
rect 454 -1281 461 -1263
rect 453 -1286 461 -1281
rect 454 -1290 461 -1286
rect 1308 -1364 1318 -1358
rect 1358 -1363 1368 -1357
rect 1408 -1363 1418 -1357
rect 1455 -1363 1465 -1357
rect 3193 -1467 3200 -1457
rect 3215 -1525 3233 -1521
rect 456 -1568 463 -1558
rect 1785 -1577 1788 -1572
rect 1823 -1577 1826 -1572
rect 1867 -1577 1870 -1572
rect 1905 -1577 1908 -1572
rect 1951 -1575 1954 -1570
rect 3209 -1579 3214 -1553
rect 3232 -1556 3239 -1538
rect 3231 -1561 3239 -1556
rect 3232 -1565 3239 -1561
rect 478 -1626 496 -1622
rect 1251 -1639 1255 -1634
rect 1279 -1639 1283 -1634
rect 1306 -1639 1310 -1634
rect 1345 -1639 1349 -1634
rect 1373 -1639 1377 -1634
rect 1400 -1639 1404 -1634
rect 1440 -1638 1444 -1633
rect 1468 -1638 1472 -1633
rect 1495 -1638 1499 -1633
rect 1531 -1638 1535 -1633
rect 472 -1680 477 -1654
rect 495 -1657 502 -1639
rect 494 -1662 502 -1657
rect 495 -1666 502 -1662
rect 481 -1877 488 -1867
rect 3213 -1884 3220 -1874
rect 503 -1935 521 -1931
rect 3235 -1942 3253 -1938
rect 497 -1989 502 -1963
rect 520 -1966 527 -1948
rect 519 -1971 527 -1966
rect 520 -1975 527 -1971
rect 3229 -1996 3234 -1970
rect 3252 -1973 3259 -1955
rect 3251 -1978 3259 -1973
rect 3252 -1982 3259 -1978
rect 477 -2232 484 -2222
rect 3262 -2270 3269 -2260
rect 499 -2290 517 -2286
rect 493 -2344 498 -2318
rect 516 -2321 523 -2303
rect 515 -2326 523 -2321
rect 516 -2330 523 -2326
rect 3284 -2328 3302 -2324
rect 3278 -2382 3283 -2356
rect 3301 -2359 3308 -2341
rect 3300 -2364 3308 -2359
rect 3301 -2368 3308 -2364
<< labels >>
rlabel metal1 1255 -1523 1259 -1519 1 pdr1
rlabel metal2 1251 -1639 1255 -1634 2 prop_1
rlabel metal1 1263 -1633 1267 -1628 1 prop1_car0
rlabel metal1 1283 -1524 1287 -1519 1 prop1_car0
rlabel metal2 1279 -1639 1283 -1634 1 carry_0
rlabel metal1 1291 -1633 1295 -1628 1 clock_car0
rlabel metal1 1310 -1524 1314 -1519 1 clock_car0
rlabel metal2 1306 -1639 1310 -1634 1 clock_in
rlabel metal1 1318 -1633 1322 -1628 1 gnd!
rlabel metal1 1349 -1524 1353 -1519 1 pdr2
rlabel metal2 1345 -1639 1349 -1634 1 prop_2
rlabel metal1 1357 -1633 1361 -1628 1 pdr1
rlabel metal1 1377 -1524 1381 -1519 1 pdr1
rlabel metal2 1373 -1639 1377 -1634 1 gen_1
rlabel metal1 1385 -1633 1389 -1628 1 clock_car0
rlabel metal1 1404 -1524 1408 -1519 1 pdr3
rlabel metal2 1400 -1639 1404 -1634 1 prop_3
rlabel metal1 1412 -1633 1416 -1628 1 pdr2
rlabel metal1 1444 -1523 1448 -1518 1 pdr2
rlabel metal2 1440 -1638 1444 -1633 1 gen_2
rlabel metal1 1452 -1632 1456 -1627 1 clock_car0
rlabel metal1 1472 -1523 1476 -1518 1 pdr4
rlabel metal2 1468 -1638 1472 -1633 1 prop_4
rlabel metal1 1480 -1632 1484 -1627 1 pdr3
rlabel metal1 1499 -1523 1503 -1518 1 pdr3
rlabel metal2 1495 -1638 1499 -1633 1 gen_3
rlabel metal1 1507 -1632 1511 -1627 1 clock_car0
rlabel metal1 1535 -1523 1539 -1518 1 pdr4
rlabel metal2 1531 -1638 1535 -1633 1 gen_4
rlabel metal1 1543 -1632 1547 -1627 7 clock_car0
rlabel metal1 1319 -1276 1323 -1271 5 vdd!
rlabel metal1 1369 -1275 1373 -1270 5 vdd!
rlabel metal1 1419 -1275 1423 -1270 5 vdd!
rlabel metal1 1466 -1275 1470 -1270 5 vdd!
rlabel metal2 1308 -1364 1314 -1358 2 clock_in
rlabel metal2 1358 -1363 1364 -1357 1 clock_in
rlabel metal2 1408 -1363 1414 -1357 1 clock_in
rlabel metal2 1455 -1363 1460 -1357 1 clock_in
rlabel metal1 1327 -1355 1331 -1350 1 pdr1
rlabel metal1 1377 -1354 1381 -1350 1 pdr2
rlabel metal1 1427 -1354 1431 -1350 1 pdr3
rlabel metal1 1474 -1354 1478 -1350 1 pdr4
rlabel metal1 1913 -1613 1917 -1609 1 gnd!
rlabel metal1 1909 -1509 1914 -1505 5 vdd!
rlabel metal2 1785 -1577 1788 -1572 1 pdr1
rlabel metal2 1823 -1577 1826 -1572 1 pdr2
rlabel metal2 1867 -1577 1870 -1572 1 pdr3
rlabel metal2 1905 -1577 1908 -1572 1 pdr4
rlabel metal1 1796 -1577 1800 -1572 1 c1
rlabel metal1 1834 -1577 1838 -1572 1 c2
rlabel metal1 1878 -1577 1882 -1572 1 c3
rlabel metal1 1916 -1577 1920 -1572 1 c4
rlabel metal1 1959 -1611 1963 -1607 1 gnd!
rlabel metal1 1955 -1507 1960 -1503 5 vdd!
rlabel metal2 1951 -1575 1954 -1570 1 clk_org
rlabel metal1 1962 -1575 1966 -1570 1 clock_in
rlabel metal1 1788 -1509 1792 -1505 5 vdd!
rlabel metal1 1826 -1509 1830 -1505 5 vdd!
rlabel metal1 1870 -1509 1874 -1505 5 vdd!
rlabel metal1 1874 -1613 1878 -1609 1 gnd!
rlabel metal1 1837 -1613 1841 -1609 1 gnd!
rlabel metal1 1797 -1613 1801 -1609 1 gnd!
rlabel metal1 118 -1387 118 -1387 5 vdd
rlabel metal1 119 -1474 119 -1474 1 gnd
rlabel metal1 151 -1456 151 -1456 1 gnd
rlabel metal1 148 -1399 148 -1399 5 vdd
rlabel metal1 120 -1737 120 -1737 5 vdd
rlabel metal1 121 -1824 121 -1824 1 gnd
rlabel metal1 153 -1806 153 -1806 1 gnd
rlabel metal1 150 -1749 150 -1749 5 vdd
rlabel metal1 128 -2029 128 -2029 5 vdd
rlabel metal1 129 -2116 129 -2116 1 gnd
rlabel metal1 161 -2098 161 -2098 1 gnd
rlabel metal1 158 -2041 158 -2041 5 vdd
rlabel metal1 116 -2395 116 -2395 5 vdd
rlabel metal1 117 -2482 117 -2482 1 gnd
rlabel metal1 149 -2464 149 -2464 1 gnd
rlabel metal1 146 -2407 146 -2407 5 vdd
rlabel metal1 103 -1436 103 -1436 3 q_a1
rlabel metal1 105 -1443 105 -1443 3 q_b1
rlabel metal1 167 -1436 167 -1436 1 gen_1
rlabel metal1 106 -1787 106 -1787 1 q_a2
rlabel metal1 106 -1794 106 -1794 1 q_b2
rlabel metal1 169 -1785 169 -1785 1 gen_2
rlabel metal1 113 -2079 113 -2079 1 q_b3
rlabel metal1 115 -2086 115 -2086 1 q_a3
rlabel metal1 176 -2077 176 -2077 1 gen_3
rlabel metal1 101 -2444 101 -2444 3 q_a4
rlabel metal1 101 -2450 101 -2450 3 q_b4
rlabel metal1 164 -2443 164 -2443 1 gen_4
rlabel metal2 457 -1287 457 -1287 1 bbar
rlabel metal1 392 -1195 392 -1195 1 vdd
rlabel metal1 393 -1275 393 -1275 1 gnd
rlabel metal1 418 -1171 418 -1171 5 vdd
rlabel metal1 392 -1273 392 -1273 1 gnd
rlabel metal1 391 -1195 391 -1195 5 vdd
rlabel metal1 374 -1249 374 -1249 1 invi
rlabel metal1 410 -1250 410 -1250 1 invo
rlabel metal2 498 -1663 498 -1663 1 bbar
rlabel metal1 433 -1571 433 -1571 1 vdd
rlabel metal1 434 -1651 434 -1651 1 gnd
rlabel metal1 459 -1547 459 -1547 5 vdd
rlabel metal1 433 -1649 433 -1649 1 gnd
rlabel metal1 432 -1571 432 -1571 5 vdd
rlabel metal1 415 -1625 415 -1625 1 invi
rlabel metal1 451 -1626 451 -1626 1 invo
rlabel metal2 523 -1972 523 -1972 1 bbar
rlabel metal1 458 -1880 458 -1880 1 vdd
rlabel metal1 459 -1960 459 -1960 1 gnd
rlabel metal1 484 -1856 484 -1856 5 vdd
rlabel metal1 458 -1958 458 -1958 1 gnd
rlabel metal1 457 -1880 457 -1880 5 vdd
rlabel metal1 440 -1934 440 -1934 1 invi
rlabel metal1 476 -1935 476 -1935 1 invo
rlabel metal2 519 -2327 519 -2327 1 bbar
rlabel metal1 454 -2235 454 -2235 1 vdd
rlabel metal1 455 -2315 455 -2315 1 gnd
rlabel metal1 480 -2211 480 -2211 5 vdd
rlabel metal1 454 -2313 454 -2313 1 gnd
rlabel metal1 453 -2235 453 -2235 5 vdd
rlabel metal1 436 -2289 436 -2289 1 invi
rlabel metal1 472 -2290 472 -2290 1 invo
rlabel metal2 3179 -1141 3179 -1141 1 bbar
rlabel metal1 3114 -1049 3114 -1049 1 vdd
rlabel metal1 3115 -1129 3115 -1129 1 gnd
rlabel metal1 3140 -1025 3140 -1025 5 vdd
rlabel metal1 3114 -1127 3114 -1127 1 gnd
rlabel metal1 3113 -1049 3113 -1049 5 vdd
rlabel metal1 3096 -1103 3096 -1103 1 invi
rlabel metal1 3132 -1104 3132 -1104 1 invo
rlabel metal2 3235 -1562 3235 -1562 1 bbar
rlabel metal1 3170 -1470 3170 -1470 1 vdd
rlabel metal1 3171 -1550 3171 -1550 1 gnd
rlabel metal1 3196 -1446 3196 -1446 5 vdd
rlabel metal1 3170 -1548 3170 -1548 1 gnd
rlabel metal1 3169 -1470 3169 -1470 5 vdd
rlabel metal1 3152 -1524 3152 -1524 1 invi
rlabel metal1 3188 -1525 3188 -1525 1 invo
rlabel metal2 3255 -1979 3255 -1979 1 bbar
rlabel metal1 3190 -1887 3190 -1887 1 vdd
rlabel metal1 3191 -1967 3191 -1967 1 gnd
rlabel metal1 3216 -1863 3216 -1863 5 vdd
rlabel metal1 3190 -1965 3190 -1965 1 gnd
rlabel metal1 3189 -1887 3189 -1887 5 vdd
rlabel metal1 3172 -1941 3172 -1941 1 invi
rlabel metal1 3208 -1942 3208 -1942 1 invo
rlabel metal2 3304 -2365 3304 -2365 1 bbar
rlabel metal1 3239 -2273 3239 -2273 1 vdd
rlabel metal1 3240 -2353 3240 -2353 1 gnd
rlabel metal1 3265 -2249 3265 -2249 5 vdd
rlabel metal1 3239 -2351 3239 -2351 1 gnd
rlabel metal1 3238 -2273 3238 -2273 5 vdd
rlabel metal1 3221 -2327 3221 -2327 1 invi
rlabel metal1 3257 -2328 3257 -2328 1 invo
rlabel metal1 433 -1242 433 -1242 1 q_a1
rlabel metal1 454 -1173 454 -1173 1 q_b1
rlabel metal1 494 -1249 494 -1249 1 prop_1
rlabel metal1 495 -1551 495 -1551 1 q_b2
rlabel metal1 474 -1619 474 -1619 1 q_a2
rlabel metal1 535 -1624 535 -1624 1 prop_2
rlabel metal1 500 -1928 500 -1928 1 q_a3
rlabel metal1 518 -1858 518 -1858 1 q_b3
rlabel metal1 561 -1933 561 -1933 1 prop_3
rlabel metal1 515 -2213 515 -2213 1 q_a4
rlabel metal1 496 -2283 496 -2283 1 q_b4
rlabel metal1 556 -2289 556 -2289 1 prop_4
rlabel metal1 3231 -1449 3231 -1449 1 carry_0
rlabel metal1 3212 -1518 3212 -1518 1 prop_1
rlabel metal1 3273 -1524 3273 -1524 1 s1
rlabel metal1 3293 -1940 3293 -1940 1 s2
rlabel metal1 3343 -2326 3343 -2326 7 s3
rlabel metal1 3219 -1102 3219 -1102 1 s4
rlabel metal1 3175 -1026 3175 -1026 5 c3
rlabel metal1 3155 -1108 3155 -1108 1 prop_4
rlabel metal1 3251 -1864 3251 -1864 1 c1
rlabel metal1 3232 -1946 3232 -1946 1 prop_1
rlabel metal1 3299 -2251 3299 -2251 1 c2
rlabel metal1 3281 -2331 3281 -2331 1 prop_3
<< end >>
