magic
tech scmos
timestamp 1731935527
<< nwell >>
rect 0 0 24 62
<< ptransistor >>
rect 11 6 13 56
<< pdiffusion >>
rect 10 6 11 56
rect 13 6 14 56
<< pdcontact >>
rect 6 6 10 56
rect 14 6 18 56
<< nsubstratencontact >>
rect 1 62 5 66
<< polysilicon >>
rect 11 56 13 59
rect 11 -9 13 6
<< metal1 >>
rect 6 66 10 69
rect 0 62 1 66
rect 5 62 10 66
rect 6 56 10 62
rect 15 -4 18 6
<< pm12contact >>
rect 6 -9 11 -4
<< metal2 >>
rect 3 -9 6 -4
<< end >>
