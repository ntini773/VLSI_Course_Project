magic
tech scmos
timestamp 1732102597
<< nwell >>
rect 3861 1452 3885 1476
rect 3900 1466 3934 1472
rect 3900 1436 3962 1466
rect 3928 1430 3962 1436
rect 3861 1397 3885 1421
rect 3878 1182 3914 1210
rect 3872 1176 3914 1182
rect 3872 1148 3908 1176
rect 4047 1134 4083 1162
rect 3868 1109 3892 1133
rect 3923 1109 3947 1133
rect 4041 1128 4083 1134
rect 4041 1100 4077 1128
rect 3496 1057 3520 1081
rect 3535 1071 3569 1077
rect 3535 1041 3597 1071
rect 4037 1061 4061 1085
rect 4092 1061 4116 1085
rect 3563 1035 3597 1041
rect 3496 1002 3520 1026
rect 4230 976 4266 1004
rect 4224 970 4266 976
rect 3497 925 3521 949
rect 3536 939 3570 945
rect 4224 942 4260 970
rect 3536 909 3598 939
rect 3564 903 3598 909
rect 3497 870 3521 894
rect 3841 887 3893 911
rect 4220 903 4244 927
rect 4275 903 4299 927
rect 4008 844 4060 868
rect 4190 837 4242 861
rect 3500 781 3524 805
rect 3539 795 3573 801
rect 3539 765 3601 795
rect 3567 759 3601 765
rect 3500 726 3524 750
rect 4476 713 4500 765
rect 4347 682 4409 706
rect 3507 656 3531 680
rect 3546 670 3580 676
rect 3546 640 3608 670
rect 3574 634 3608 640
rect 3507 601 3531 625
rect 3803 620 3865 644
rect 3977 643 4039 667
rect 4151 647 4213 671
rect 3529 423 3565 463
rect 3571 416 3595 456
rect 3529 314 3565 354
rect 3571 307 3595 347
rect 3875 328 3927 352
rect 3684 299 3721 325
rect 3684 254 3721 280
rect 3530 195 3566 235
rect 3572 188 3596 228
rect 3684 210 3721 236
rect 3684 172 3721 204
rect 3534 87 3570 127
rect 3576 80 3600 120
<< ntransistor >>
rect 3872 1438 3874 1444
rect 3911 1389 3913 1401
rect 3921 1389 3923 1401
rect 3939 1389 3941 1401
rect 3949 1389 3951 1401
rect 3872 1383 3874 1389
rect 3943 1197 3955 1199
rect 3943 1187 3955 1189
rect 3943 1169 3955 1171
rect 3943 1159 3955 1161
rect 4112 1149 4124 1151
rect 4112 1139 4124 1141
rect 3900 1120 3906 1122
rect 3955 1120 3961 1122
rect 4112 1121 4124 1123
rect 4112 1111 4124 1113
rect 4069 1072 4075 1074
rect 4124 1072 4130 1074
rect 3507 1043 3509 1049
rect 3546 994 3548 1006
rect 3556 994 3558 1006
rect 3574 994 3576 1006
rect 3584 994 3586 1006
rect 3507 988 3509 994
rect 4295 991 4307 993
rect 4295 981 4307 983
rect 4295 963 4307 965
rect 4295 953 4307 955
rect 3508 911 3510 917
rect 4252 914 4258 916
rect 4307 914 4313 916
rect 3905 898 3925 900
rect 3547 862 3549 874
rect 3557 862 3559 874
rect 3575 862 3577 874
rect 3585 862 3587 874
rect 3508 856 3510 862
rect 4072 855 4092 857
rect 4254 848 4274 850
rect 3511 767 3513 773
rect 3550 718 3552 730
rect 3560 718 3562 730
rect 3578 718 3580 730
rect 3588 718 3590 730
rect 3511 712 3513 718
rect 4487 681 4489 701
rect 3518 642 3520 648
rect 4329 608 4429 610
rect 3557 593 3559 605
rect 3567 593 3569 605
rect 3585 593 3587 605
rect 3595 593 3597 605
rect 4141 600 4241 602
rect 3518 587 3520 593
rect 3960 590 4060 592
rect 3792 582 3892 584
rect 4331 499 4431 501
rect 4139 489 4239 491
rect 3959 479 4059 481
rect 3540 380 3542 400
rect 3551 380 3553 400
rect 3582 398 3584 408
rect 3744 371 3746 471
rect 3791 468 3891 470
rect 3824 370 3924 372
rect 3939 339 3959 341
rect 3737 310 3747 312
rect 3540 271 3542 291
rect 3551 271 3553 291
rect 3582 289 3584 299
rect 3737 267 3747 269
rect 3737 259 3747 261
rect 3737 223 3747 225
rect 3737 215 3747 217
rect 3541 152 3543 172
rect 3552 152 3554 172
rect 3583 170 3585 180
rect 3737 179 3747 181
rect 3545 44 3547 64
rect 3556 44 3558 64
rect 3587 62 3589 72
<< ptransistor >>
rect 3872 1458 3874 1470
rect 3911 1442 3913 1466
rect 3921 1442 3923 1466
rect 3939 1436 3941 1460
rect 3949 1436 3951 1460
rect 3872 1403 3874 1415
rect 3884 1197 3908 1199
rect 3884 1187 3908 1189
rect 3878 1169 3902 1171
rect 3878 1159 3902 1161
rect 4053 1149 4077 1151
rect 4053 1139 4077 1141
rect 3874 1120 3886 1122
rect 3929 1120 3941 1122
rect 4047 1121 4071 1123
rect 4047 1111 4071 1113
rect 3507 1063 3509 1075
rect 4043 1072 4055 1074
rect 4098 1072 4110 1074
rect 3546 1047 3548 1071
rect 3556 1047 3558 1071
rect 3574 1041 3576 1065
rect 3584 1041 3586 1065
rect 3507 1008 3509 1020
rect 4236 991 4260 993
rect 4236 981 4260 983
rect 4230 963 4254 965
rect 4230 953 4254 955
rect 3508 931 3510 943
rect 3547 915 3549 939
rect 3557 915 3559 939
rect 3575 909 3577 933
rect 3585 909 3587 933
rect 4226 914 4238 916
rect 4281 914 4293 916
rect 3508 876 3510 888
rect 3847 898 3887 900
rect 4014 855 4054 857
rect 4196 848 4236 850
rect 3511 787 3513 799
rect 3550 771 3552 795
rect 3560 771 3562 795
rect 3578 765 3580 789
rect 3588 765 3590 789
rect 3511 732 3513 744
rect 4487 719 4489 759
rect 4353 693 4403 695
rect 3518 662 3520 674
rect 3557 646 3559 670
rect 3567 646 3569 670
rect 3585 640 3587 664
rect 3595 640 3597 664
rect 4157 658 4207 660
rect 3983 654 4033 656
rect 3518 607 3520 619
rect 3809 631 3859 633
rect 3540 429 3542 449
rect 3551 429 3553 449
rect 3582 422 3584 442
rect 3540 320 3542 340
rect 3551 320 3553 340
rect 3881 339 3921 341
rect 3582 313 3584 333
rect 3690 310 3715 312
rect 3690 265 3715 267
rect 3690 221 3715 223
rect 3541 201 3543 221
rect 3552 201 3554 221
rect 3583 194 3585 214
rect 3690 191 3715 193
rect 3690 183 3715 185
rect 3545 93 3547 113
rect 3556 93 3558 113
rect 3587 86 3589 106
<< ndiffusion >>
rect 3871 1438 3872 1444
rect 3874 1438 3875 1444
rect 3910 1389 3911 1401
rect 3913 1389 3921 1401
rect 3923 1389 3924 1401
rect 3938 1389 3939 1401
rect 3941 1389 3949 1401
rect 3951 1389 3952 1401
rect 3871 1383 3872 1389
rect 3874 1383 3875 1389
rect 3943 1199 3955 1200
rect 3943 1189 3955 1197
rect 3943 1186 3955 1187
rect 3943 1171 3955 1172
rect 3943 1161 3955 1169
rect 3943 1158 3955 1159
rect 4112 1151 4124 1152
rect 4112 1141 4124 1149
rect 4112 1138 4124 1139
rect 3900 1122 3906 1123
rect 4112 1123 4124 1124
rect 3955 1122 3961 1123
rect 3900 1119 3906 1120
rect 3955 1119 3961 1120
rect 4112 1113 4124 1121
rect 4112 1110 4124 1111
rect 4069 1074 4075 1075
rect 4124 1074 4130 1075
rect 3506 1043 3507 1049
rect 3509 1043 3510 1049
rect 4069 1071 4075 1072
rect 4124 1071 4130 1072
rect 3545 994 3546 1006
rect 3548 994 3556 1006
rect 3558 994 3559 1006
rect 3573 994 3574 1006
rect 3576 994 3584 1006
rect 3586 994 3587 1006
rect 3506 988 3507 994
rect 3509 988 3510 994
rect 4295 993 4307 994
rect 4295 983 4307 991
rect 4295 980 4307 981
rect 4295 965 4307 966
rect 4295 955 4307 963
rect 4295 952 4307 953
rect 3507 911 3508 917
rect 3510 911 3511 917
rect 4252 916 4258 917
rect 4307 916 4313 917
rect 4252 913 4258 914
rect 4307 913 4313 914
rect 3905 900 3925 901
rect 3905 897 3925 898
rect 3546 862 3547 874
rect 3549 862 3557 874
rect 3559 862 3560 874
rect 3574 862 3575 874
rect 3577 862 3585 874
rect 3587 862 3588 874
rect 3507 856 3508 862
rect 3510 856 3511 862
rect 4072 857 4092 858
rect 4072 854 4092 855
rect 4254 850 4274 851
rect 4254 847 4274 848
rect 3510 767 3511 773
rect 3513 767 3514 773
rect 3549 718 3550 730
rect 3552 718 3560 730
rect 3562 718 3563 730
rect 3577 718 3578 730
rect 3580 718 3588 730
rect 3590 718 3591 730
rect 3510 712 3511 718
rect 3513 712 3514 718
rect 4486 681 4487 701
rect 4489 681 4490 701
rect 3517 642 3518 648
rect 3520 642 3521 648
rect 4329 610 4429 611
rect 4329 607 4429 608
rect 3556 593 3557 605
rect 3559 593 3567 605
rect 3569 593 3570 605
rect 3584 593 3585 605
rect 3587 593 3595 605
rect 3597 593 3598 605
rect 4141 602 4241 603
rect 4141 599 4241 600
rect 3517 587 3518 593
rect 3520 587 3521 593
rect 3960 592 4060 593
rect 3960 589 4060 590
rect 3792 584 3892 585
rect 3792 581 3892 582
rect 4331 501 4431 502
rect 4331 498 4431 499
rect 4139 491 4239 492
rect 4139 488 4239 489
rect 3959 481 4059 482
rect 3959 478 4059 479
rect 3539 380 3540 400
rect 3542 380 3551 400
rect 3553 380 3554 400
rect 3581 398 3582 408
rect 3584 398 3585 408
rect 3743 371 3744 471
rect 3746 371 3747 471
rect 3791 470 3891 471
rect 3791 467 3891 468
rect 3824 372 3924 373
rect 3824 369 3924 370
rect 3939 341 3959 342
rect 3939 338 3959 339
rect 3737 312 3747 313
rect 3737 309 3747 310
rect 3539 271 3540 291
rect 3542 271 3551 291
rect 3553 271 3554 291
rect 3581 289 3582 299
rect 3584 289 3585 299
rect 3737 269 3747 270
rect 3737 266 3747 267
rect 3737 261 3747 262
rect 3737 258 3747 259
rect 3737 225 3747 226
rect 3737 222 3747 223
rect 3737 217 3747 218
rect 3737 214 3747 215
rect 3540 152 3541 172
rect 3543 152 3552 172
rect 3554 152 3555 172
rect 3582 170 3583 180
rect 3585 170 3586 180
rect 3737 181 3747 182
rect 3737 178 3747 179
rect 3544 44 3545 64
rect 3547 44 3556 64
rect 3558 44 3559 64
rect 3586 62 3587 72
rect 3589 62 3590 72
<< pdiffusion >>
rect 3871 1458 3872 1470
rect 3874 1458 3875 1470
rect 3910 1442 3911 1466
rect 3913 1442 3915 1466
rect 3919 1442 3921 1466
rect 3923 1442 3924 1466
rect 3938 1436 3939 1460
rect 3941 1436 3943 1460
rect 3947 1436 3949 1460
rect 3951 1436 3952 1460
rect 3871 1403 3872 1415
rect 3874 1403 3875 1415
rect 3884 1199 3908 1200
rect 3884 1195 3908 1197
rect 3884 1189 3908 1191
rect 3884 1186 3908 1187
rect 3878 1171 3902 1172
rect 3878 1167 3902 1169
rect 3878 1161 3902 1163
rect 3878 1158 3902 1159
rect 4053 1151 4077 1152
rect 4053 1147 4077 1149
rect 4053 1141 4077 1143
rect 4053 1138 4077 1139
rect 3874 1122 3886 1123
rect 3929 1122 3941 1123
rect 4047 1123 4071 1124
rect 3874 1119 3886 1120
rect 3929 1119 3941 1120
rect 4047 1119 4071 1121
rect 4047 1113 4071 1115
rect 4047 1110 4071 1111
rect 3506 1063 3507 1075
rect 3509 1063 3510 1075
rect 4043 1074 4055 1075
rect 4098 1074 4110 1075
rect 4043 1071 4055 1072
rect 3545 1047 3546 1071
rect 3548 1047 3550 1071
rect 3554 1047 3556 1071
rect 3558 1047 3559 1071
rect 4098 1071 4110 1072
rect 3573 1041 3574 1065
rect 3576 1041 3578 1065
rect 3582 1041 3584 1065
rect 3586 1041 3587 1065
rect 3506 1008 3507 1020
rect 3509 1008 3510 1020
rect 4236 993 4260 994
rect 4236 989 4260 991
rect 4236 983 4260 985
rect 4236 980 4260 981
rect 4230 965 4254 966
rect 4230 961 4254 963
rect 4230 955 4254 957
rect 4230 952 4254 953
rect 3507 931 3508 943
rect 3510 931 3511 943
rect 3546 915 3547 939
rect 3549 915 3551 939
rect 3555 915 3557 939
rect 3559 915 3560 939
rect 3574 909 3575 933
rect 3577 909 3579 933
rect 3583 909 3585 933
rect 3587 909 3588 933
rect 4226 916 4238 917
rect 4281 916 4293 917
rect 4226 913 4238 914
rect 4281 913 4293 914
rect 3507 876 3508 888
rect 3510 876 3511 888
rect 3847 900 3887 901
rect 3847 897 3887 898
rect 4014 857 4054 858
rect 4014 854 4054 855
rect 4196 850 4236 851
rect 4196 847 4236 848
rect 3510 787 3511 799
rect 3513 787 3514 799
rect 3549 771 3550 795
rect 3552 771 3554 795
rect 3558 771 3560 795
rect 3562 771 3563 795
rect 3577 765 3578 789
rect 3580 765 3582 789
rect 3586 765 3588 789
rect 3590 765 3591 789
rect 3510 732 3511 744
rect 3513 732 3514 744
rect 4486 719 4487 759
rect 4489 719 4490 759
rect 4353 695 4403 696
rect 4353 692 4403 693
rect 3517 662 3518 674
rect 3520 662 3521 674
rect 3556 646 3557 670
rect 3559 646 3561 670
rect 3565 646 3567 670
rect 3569 646 3570 670
rect 3584 640 3585 664
rect 3587 640 3589 664
rect 3593 640 3595 664
rect 3597 640 3598 664
rect 3983 656 4033 657
rect 4157 660 4207 661
rect 4157 657 4207 658
rect 3983 653 4033 654
rect 3517 607 3518 619
rect 3520 607 3521 619
rect 3809 633 3859 634
rect 3809 630 3859 631
rect 3539 429 3540 449
rect 3542 429 3546 449
rect 3550 429 3551 449
rect 3553 429 3554 449
rect 3581 422 3582 442
rect 3584 422 3585 442
rect 3881 341 3921 342
rect 3539 320 3540 340
rect 3542 320 3546 340
rect 3550 320 3551 340
rect 3553 320 3554 340
rect 3881 338 3921 339
rect 3581 313 3582 333
rect 3584 313 3585 333
rect 3690 312 3715 313
rect 3690 309 3715 310
rect 3690 267 3715 268
rect 3690 264 3715 265
rect 3690 223 3715 224
rect 3540 201 3541 221
rect 3543 201 3547 221
rect 3551 201 3552 221
rect 3554 201 3555 221
rect 3690 220 3715 221
rect 3582 194 3583 214
rect 3585 194 3586 214
rect 3690 193 3715 194
rect 3690 190 3715 191
rect 3690 185 3715 186
rect 3690 182 3715 183
rect 3544 93 3545 113
rect 3547 93 3551 113
rect 3555 93 3556 113
rect 3558 93 3559 113
rect 3586 86 3587 106
rect 3589 86 3590 106
<< ndcontact >>
rect 3867 1438 3871 1444
rect 3875 1438 3879 1444
rect 3906 1389 3910 1401
rect 3924 1389 3928 1401
rect 3934 1389 3938 1401
rect 3952 1389 3956 1401
rect 3867 1383 3871 1389
rect 3875 1383 3879 1389
rect 3943 1200 3955 1204
rect 3943 1182 3955 1186
rect 3943 1172 3955 1176
rect 3943 1154 3955 1158
rect 4112 1152 4124 1156
rect 4112 1134 4124 1138
rect 3900 1123 3906 1127
rect 3955 1123 3961 1127
rect 4112 1124 4124 1128
rect 3900 1115 3906 1119
rect 3955 1115 3961 1119
rect 4112 1106 4124 1110
rect 4069 1075 4075 1079
rect 4124 1075 4130 1079
rect 3502 1043 3506 1049
rect 3510 1043 3514 1049
rect 4069 1067 4075 1071
rect 4124 1067 4130 1071
rect 3541 994 3545 1006
rect 3559 994 3563 1006
rect 3569 994 3573 1006
rect 3587 994 3591 1006
rect 4295 994 4307 998
rect 3502 988 3506 994
rect 3510 988 3514 994
rect 4295 976 4307 980
rect 4295 966 4307 970
rect 4295 948 4307 952
rect 3503 911 3507 917
rect 3511 911 3515 917
rect 4252 917 4258 921
rect 4307 917 4313 921
rect 4252 909 4258 913
rect 4307 909 4313 913
rect 3905 901 3925 905
rect 3905 893 3925 897
rect 3542 862 3546 874
rect 3560 862 3564 874
rect 3570 862 3574 874
rect 3588 862 3592 874
rect 3503 856 3507 862
rect 3511 856 3515 862
rect 4072 858 4092 862
rect 4072 850 4092 854
rect 4254 851 4274 855
rect 4254 843 4274 847
rect 3506 767 3510 773
rect 3514 767 3518 773
rect 3545 718 3549 730
rect 3563 718 3567 730
rect 3573 718 3577 730
rect 3591 718 3595 730
rect 3506 712 3510 718
rect 3514 712 3518 718
rect 4482 681 4486 701
rect 4490 681 4494 701
rect 3513 642 3517 648
rect 3521 642 3525 648
rect 4329 611 4429 615
rect 3552 593 3556 605
rect 3570 593 3574 605
rect 3580 593 3584 605
rect 3598 593 3602 605
rect 4141 603 4241 607
rect 4329 603 4429 607
rect 3513 587 3517 593
rect 3521 587 3525 593
rect 3960 593 4060 597
rect 4141 595 4241 599
rect 3792 585 3892 589
rect 3960 585 4060 589
rect 3792 577 3892 581
rect 4331 502 4431 506
rect 4139 492 4239 496
rect 4331 494 4431 498
rect 3959 482 4059 486
rect 4139 484 4239 488
rect 3535 380 3539 400
rect 3554 380 3558 400
rect 3577 398 3581 408
rect 3585 398 3589 408
rect 3739 371 3743 471
rect 3747 371 3751 471
rect 3791 471 3891 475
rect 3959 474 4059 478
rect 3791 463 3891 467
rect 3824 373 3924 377
rect 3824 365 3924 369
rect 3939 342 3959 346
rect 3939 334 3959 338
rect 3737 313 3747 317
rect 3737 305 3747 309
rect 3535 271 3539 291
rect 3554 271 3558 291
rect 3577 289 3581 299
rect 3585 289 3589 299
rect 3737 270 3747 274
rect 3737 262 3747 266
rect 3737 254 3747 258
rect 3737 226 3747 230
rect 3737 218 3747 222
rect 3737 210 3747 214
rect 3536 152 3540 172
rect 3555 152 3559 172
rect 3578 170 3582 180
rect 3586 170 3590 180
rect 3737 182 3747 186
rect 3737 174 3747 178
rect 3540 44 3544 64
rect 3559 44 3563 64
rect 3582 62 3586 72
rect 3590 62 3594 72
<< pdcontact >>
rect 3867 1458 3871 1470
rect 3875 1458 3879 1470
rect 3906 1442 3910 1466
rect 3915 1442 3919 1466
rect 3924 1442 3928 1466
rect 3934 1436 3938 1460
rect 3943 1436 3947 1460
rect 3952 1436 3956 1460
rect 3867 1403 3871 1415
rect 3875 1403 3879 1415
rect 3884 1200 3908 1204
rect 3884 1191 3908 1195
rect 3884 1182 3908 1186
rect 3878 1172 3902 1176
rect 3878 1163 3902 1167
rect 3878 1154 3902 1158
rect 4053 1152 4077 1156
rect 4053 1143 4077 1147
rect 4053 1134 4077 1138
rect 3874 1123 3886 1127
rect 3929 1123 3941 1127
rect 4047 1124 4071 1128
rect 3874 1115 3886 1119
rect 3929 1115 3941 1119
rect 4047 1115 4071 1119
rect 4047 1106 4071 1110
rect 4043 1075 4055 1079
rect 3502 1063 3506 1075
rect 3510 1063 3514 1075
rect 4098 1075 4110 1079
rect 3541 1047 3545 1071
rect 3550 1047 3554 1071
rect 3559 1047 3563 1071
rect 4043 1067 4055 1071
rect 4098 1067 4110 1071
rect 3569 1041 3573 1065
rect 3578 1041 3582 1065
rect 3587 1041 3591 1065
rect 3502 1008 3506 1020
rect 3510 1008 3514 1020
rect 4236 994 4260 998
rect 4236 985 4260 989
rect 4236 976 4260 980
rect 4230 966 4254 970
rect 4230 957 4254 961
rect 4230 948 4254 952
rect 3503 931 3507 943
rect 3511 931 3515 943
rect 3542 915 3546 939
rect 3551 915 3555 939
rect 3560 915 3564 939
rect 3570 909 3574 933
rect 3579 909 3583 933
rect 3588 909 3592 933
rect 4226 917 4238 921
rect 4281 917 4293 921
rect 4226 909 4238 913
rect 4281 909 4293 913
rect 3503 876 3507 888
rect 3511 876 3515 888
rect 3847 901 3887 905
rect 3847 893 3887 897
rect 4014 858 4054 862
rect 4014 850 4054 854
rect 4196 851 4236 855
rect 4196 843 4236 847
rect 3506 787 3510 799
rect 3514 787 3518 799
rect 3545 771 3549 795
rect 3554 771 3558 795
rect 3563 771 3567 795
rect 3573 765 3577 789
rect 3582 765 3586 789
rect 3591 765 3595 789
rect 3506 732 3510 744
rect 3514 732 3518 744
rect 4482 719 4486 759
rect 4490 719 4494 759
rect 4353 696 4403 700
rect 4353 688 4403 692
rect 3513 662 3517 674
rect 3521 662 3525 674
rect 3552 646 3556 670
rect 3561 646 3565 670
rect 3570 646 3574 670
rect 3580 640 3584 664
rect 3589 640 3593 664
rect 3598 640 3602 664
rect 3983 657 4033 661
rect 4157 661 4207 665
rect 4157 653 4207 657
rect 3983 649 4033 653
rect 3513 607 3517 619
rect 3521 607 3525 619
rect 3809 634 3859 638
rect 3809 626 3859 630
rect 3535 429 3539 449
rect 3546 429 3550 449
rect 3554 429 3558 449
rect 3577 422 3581 442
rect 3585 422 3589 442
rect 3881 342 3921 346
rect 3535 320 3539 340
rect 3546 320 3550 340
rect 3554 320 3558 340
rect 3881 334 3921 338
rect 3577 313 3581 333
rect 3585 313 3589 333
rect 3690 313 3715 317
rect 3690 305 3715 309
rect 3690 268 3715 272
rect 3690 260 3715 264
rect 3690 224 3715 228
rect 3536 201 3540 221
rect 3547 201 3551 221
rect 3555 201 3559 221
rect 3690 216 3715 220
rect 3578 194 3582 214
rect 3586 194 3590 214
rect 3690 194 3715 198
rect 3690 186 3715 190
rect 3690 178 3715 182
rect 3540 93 3544 113
rect 3551 93 3555 113
rect 3559 93 3563 113
rect 3582 86 3586 106
rect 3590 86 3594 106
<< psubstratepcontact >>
rect 3591 389 3596 393
rect 3591 280 3596 284
rect 3592 161 3597 165
rect 3596 53 3601 57
<< nsubstratencontact >>
rect 3837 888 3841 892
rect 4004 845 4008 849
rect 4186 838 4190 842
rect 4477 765 4481 769
rect 4342 701 4347 705
rect 4146 666 4151 670
rect 3972 662 3977 666
rect 3798 639 3803 643
rect 3535 454 3539 460
rect 3587 449 3591 453
rect 3535 345 3539 351
rect 3587 340 3591 344
rect 3871 329 3875 333
rect 3536 226 3540 232
rect 3588 221 3592 225
rect 3540 118 3544 124
rect 3592 113 3596 117
<< polysilicon >>
rect 3872 1470 3874 1473
rect 3911 1466 3913 1469
rect 3921 1466 3923 1469
rect 3872 1444 3874 1458
rect 3939 1460 3941 1463
rect 3949 1460 3951 1463
rect 3872 1435 3874 1438
rect 3911 1433 3913 1442
rect 3921 1432 3923 1442
rect 3872 1415 3874 1418
rect 3872 1389 3874 1403
rect 3911 1401 3913 1428
rect 3921 1401 3923 1427
rect 3939 1425 3941 1436
rect 3939 1401 3941 1421
rect 3949 1414 3951 1436
rect 3949 1401 3951 1410
rect 3911 1386 3913 1389
rect 3921 1386 3923 1389
rect 3939 1386 3941 1389
rect 3949 1386 3951 1389
rect 3872 1380 3874 1383
rect 3881 1197 3884 1199
rect 3908 1197 3930 1199
rect 3934 1197 3943 1199
rect 3955 1197 3958 1199
rect 3881 1187 3884 1189
rect 3908 1187 3919 1189
rect 3923 1187 3943 1189
rect 3955 1187 3958 1189
rect 3875 1169 3878 1171
rect 3902 1169 3912 1171
rect 3917 1169 3943 1171
rect 3955 1169 3958 1171
rect 3875 1159 3878 1161
rect 3902 1159 3911 1161
rect 3916 1159 3943 1161
rect 3955 1159 3958 1161
rect 4050 1149 4053 1151
rect 4077 1149 4099 1151
rect 4103 1149 4112 1151
rect 4124 1149 4127 1151
rect 4050 1139 4053 1141
rect 4077 1139 4088 1141
rect 4092 1139 4112 1141
rect 4124 1139 4127 1141
rect 3871 1120 3874 1122
rect 3886 1120 3900 1122
rect 3906 1120 3909 1122
rect 3926 1120 3929 1122
rect 3941 1120 3955 1122
rect 3961 1120 3964 1122
rect 4044 1121 4047 1123
rect 4071 1121 4081 1123
rect 4086 1121 4112 1123
rect 4124 1121 4127 1123
rect 4044 1111 4047 1113
rect 4071 1111 4080 1113
rect 4085 1111 4112 1113
rect 4124 1111 4127 1113
rect 3507 1075 3509 1078
rect 3546 1071 3548 1074
rect 3556 1071 3558 1074
rect 4040 1072 4043 1074
rect 4055 1072 4069 1074
rect 4075 1072 4078 1074
rect 4095 1072 4098 1074
rect 4110 1072 4124 1074
rect 4130 1072 4133 1074
rect 3507 1049 3509 1063
rect 3574 1065 3576 1068
rect 3584 1065 3586 1068
rect 3507 1040 3509 1043
rect 3546 1038 3548 1047
rect 3556 1037 3558 1047
rect 3507 1020 3509 1023
rect 3507 994 3509 1008
rect 3546 1006 3548 1033
rect 3556 1006 3558 1032
rect 3574 1030 3576 1041
rect 3574 1006 3576 1026
rect 3584 1019 3586 1041
rect 3584 1006 3586 1015
rect 3546 991 3548 994
rect 3556 991 3558 994
rect 3574 991 3576 994
rect 3584 991 3586 994
rect 4233 991 4236 993
rect 4260 991 4282 993
rect 4286 991 4295 993
rect 4307 991 4310 993
rect 3507 985 3509 988
rect 4233 981 4236 983
rect 4260 981 4271 983
rect 4275 981 4295 983
rect 4307 981 4310 983
rect 4227 963 4230 965
rect 4254 963 4264 965
rect 4269 963 4295 965
rect 4307 963 4310 965
rect 4227 953 4230 955
rect 4254 953 4263 955
rect 4268 953 4295 955
rect 4307 953 4310 955
rect 3508 943 3510 946
rect 3547 939 3549 942
rect 3557 939 3559 942
rect 3508 917 3510 931
rect 3575 933 3577 936
rect 3585 933 3587 936
rect 3508 908 3510 911
rect 3547 906 3549 915
rect 3557 905 3559 915
rect 4223 914 4226 916
rect 4238 914 4252 916
rect 4258 914 4261 916
rect 4278 914 4281 916
rect 4293 914 4307 916
rect 4313 914 4316 916
rect 3508 888 3510 891
rect 3508 862 3510 876
rect 3547 874 3549 901
rect 3557 874 3559 900
rect 3575 898 3577 909
rect 3575 874 3577 894
rect 3585 887 3587 909
rect 3844 898 3847 900
rect 3887 898 3905 900
rect 3925 898 3929 900
rect 3585 874 3587 883
rect 3547 859 3549 862
rect 3557 859 3559 862
rect 3575 859 3577 862
rect 3585 859 3587 862
rect 3508 853 3510 856
rect 4011 855 4014 857
rect 4054 855 4072 857
rect 4092 855 4096 857
rect 4193 848 4196 850
rect 4236 848 4254 850
rect 4274 848 4278 850
rect 3511 799 3513 802
rect 3550 795 3552 798
rect 3560 795 3562 798
rect 3511 773 3513 787
rect 3578 789 3580 792
rect 3588 789 3590 792
rect 3511 764 3513 767
rect 3550 762 3552 771
rect 3560 761 3562 771
rect 3511 744 3513 747
rect 3511 718 3513 732
rect 3550 730 3552 757
rect 3560 730 3562 756
rect 3578 754 3580 765
rect 3578 730 3580 750
rect 3588 743 3590 765
rect 4487 759 4489 762
rect 3588 730 3590 739
rect 3550 715 3552 718
rect 3560 715 3562 718
rect 3578 715 3580 718
rect 3588 715 3590 718
rect 3511 709 3513 712
rect 4487 701 4489 719
rect 4350 693 4353 695
rect 4403 693 4426 695
rect 4487 677 4489 681
rect 3518 674 3520 677
rect 3557 670 3559 673
rect 3567 670 3569 673
rect 3518 648 3520 662
rect 3585 664 3587 667
rect 3595 664 3597 667
rect 3518 639 3520 642
rect 3557 637 3559 646
rect 3567 636 3569 646
rect 4154 658 4157 660
rect 4207 658 4230 660
rect 3980 654 3983 656
rect 4033 654 4056 656
rect 3518 619 3520 622
rect 3518 593 3520 607
rect 3557 605 3559 632
rect 3567 605 3569 631
rect 3585 629 3587 640
rect 3585 605 3587 625
rect 3595 618 3597 640
rect 3806 631 3809 633
rect 3859 631 3882 633
rect 3595 605 3597 614
rect 4317 608 4329 610
rect 4429 608 4432 610
rect 4129 600 4141 602
rect 4241 600 4244 602
rect 3557 590 3559 593
rect 3567 590 3569 593
rect 3585 590 3587 593
rect 3595 590 3597 593
rect 3948 590 3960 592
rect 4060 590 4063 592
rect 3518 584 3520 587
rect 3780 582 3792 584
rect 3892 582 3895 584
rect 4319 499 4331 501
rect 4431 499 4434 501
rect 4127 489 4139 491
rect 4239 489 4242 491
rect 3947 479 3959 481
rect 4059 479 4062 481
rect 3744 471 3746 474
rect 3540 449 3542 452
rect 3551 449 3553 452
rect 3582 442 3584 446
rect 3540 400 3542 429
rect 3551 400 3553 429
rect 3582 408 3584 422
rect 3582 395 3584 398
rect 3540 377 3542 380
rect 3551 377 3553 380
rect 3779 468 3791 470
rect 3891 468 3894 470
rect 3744 359 3746 371
rect 3821 370 3824 372
rect 3924 370 3936 372
rect 3540 340 3542 343
rect 3551 340 3553 343
rect 3878 339 3881 341
rect 3921 339 3939 341
rect 3959 339 3963 341
rect 3582 333 3584 337
rect 3540 291 3542 320
rect 3551 291 3553 320
rect 3582 299 3584 313
rect 3687 310 3690 312
rect 3715 310 3737 312
rect 3747 310 3750 312
rect 3582 286 3584 289
rect 3540 268 3542 271
rect 3551 268 3553 271
rect 3728 267 3737 269
rect 3747 267 3750 269
rect 3687 265 3690 267
rect 3715 265 3725 267
rect 3723 261 3725 265
rect 3723 259 3737 261
rect 3747 259 3750 261
rect 3541 221 3543 224
rect 3552 221 3554 224
rect 3728 223 3737 225
rect 3747 223 3750 225
rect 3687 221 3690 223
rect 3715 221 3725 223
rect 3583 214 3585 218
rect 3723 217 3725 221
rect 3723 215 3737 217
rect 3747 215 3750 217
rect 3541 172 3543 201
rect 3552 172 3554 201
rect 3583 180 3585 194
rect 3687 191 3690 193
rect 3715 191 3734 193
rect 3687 183 3690 185
rect 3715 183 3726 185
rect 3722 181 3726 183
rect 3722 179 3737 181
rect 3747 179 3750 181
rect 3722 178 3726 179
rect 3583 167 3585 170
rect 3541 149 3543 152
rect 3552 149 3554 152
rect 3545 113 3547 116
rect 3556 113 3558 116
rect 3587 106 3589 110
rect 3545 64 3547 93
rect 3556 64 3558 93
rect 3587 72 3589 86
rect 3587 59 3589 62
rect 3545 41 3547 44
rect 3556 41 3558 44
<< polycontact >>
rect 3868 1447 3872 1451
rect 3868 1392 3872 1396
rect 3937 1421 3941 1425
rect 3948 1410 3952 1414
rect 3930 1196 3934 1200
rect 3919 1185 3923 1189
rect 4099 1148 4103 1152
rect 4088 1137 4092 1141
rect 3893 1116 3897 1120
rect 3948 1116 3952 1120
rect 3503 1052 3507 1056
rect 4062 1068 4066 1072
rect 4117 1068 4121 1072
rect 3503 997 3507 1001
rect 3572 1026 3576 1030
rect 3583 1015 3587 1019
rect 4282 990 4286 994
rect 4271 979 4275 983
rect 3504 920 3508 924
rect 4245 910 4249 914
rect 4300 910 4304 914
rect 3504 865 3508 869
rect 3573 894 3577 898
rect 3584 883 3588 887
rect 3507 776 3511 780
rect 3507 721 3511 725
rect 3576 750 3580 754
rect 3587 739 3591 743
rect 4482 704 4487 709
rect 3514 651 3518 655
rect 3514 596 3518 600
rect 3583 625 3587 629
rect 3594 614 3598 618
rect 3536 403 3540 407
rect 3547 410 3551 414
rect 3578 411 3582 415
rect 3536 294 3540 298
rect 3547 301 3551 305
rect 3578 302 3582 306
rect 3724 306 3729 310
rect 3730 269 3734 273
rect 3729 254 3734 259
rect 3730 225 3734 229
rect 3537 175 3541 179
rect 3548 182 3552 186
rect 3729 210 3734 215
rect 3722 198 3726 202
rect 3579 183 3583 187
rect 3730 187 3734 191
rect 3722 174 3726 178
rect 3541 67 3545 71
rect 3552 74 3556 78
rect 3583 75 3587 79
<< metal1 >>
rect 3866 1476 3894 1479
rect 3867 1470 3870 1476
rect 3891 1475 3894 1476
rect 3891 1472 3962 1475
rect 3706 1446 3853 1449
rect 3501 1081 3529 1084
rect 3502 1075 3505 1081
rect 3526 1080 3529 1081
rect 3526 1077 3597 1080
rect 3473 1051 3488 1054
rect 3493 1052 3503 1055
rect 3511 1055 3514 1063
rect 3541 1071 3544 1077
rect 3560 1071 3563 1077
rect 3511 1052 3532 1055
rect 3511 1049 3514 1052
rect 3502 1039 3505 1043
rect 3496 1037 3520 1039
rect 3496 1036 3514 1037
rect 3519 1036 3520 1037
rect 3529 1029 3532 1052
rect 3570 1071 3590 1074
rect 3570 1065 3573 1071
rect 3587 1065 3590 1071
rect 3551 1044 3554 1047
rect 3551 1041 3569 1044
rect 3579 1034 3582 1041
rect 3579 1031 3596 1034
rect 3501 1028 3520 1029
rect 3496 1026 3520 1028
rect 3529 1026 3572 1029
rect 3502 1020 3505 1026
rect 3593 1020 3596 1031
rect 3558 1015 3583 1018
rect 3593 1016 3606 1020
rect 3558 1013 3561 1015
rect 3473 997 3488 1000
rect 3493 997 3503 1000
rect 3511 1000 3514 1008
rect 3523 1010 3561 1013
rect 3593 1012 3596 1016
rect 3523 1000 3526 1010
rect 3564 1009 3596 1012
rect 3564 1006 3567 1009
rect 3511 997 3526 1000
rect 3511 994 3514 997
rect 3563 1003 3569 1006
rect 3502 984 3505 988
rect 3523 987 3528 990
rect 3541 990 3544 994
rect 3588 990 3591 994
rect 3533 987 3597 990
rect 3523 984 3526 987
rect 3496 981 3526 984
rect 3602 981 3606 1016
rect 3502 949 3530 952
rect 3503 943 3506 949
rect 3527 948 3530 949
rect 3527 945 3598 948
rect 3473 919 3489 922
rect 3494 920 3504 923
rect 3512 923 3515 931
rect 3542 939 3545 945
rect 3561 939 3564 945
rect 3512 920 3533 923
rect 3512 917 3515 920
rect 3503 907 3506 911
rect 3497 905 3521 907
rect 3497 904 3515 905
rect 3520 904 3521 905
rect 3530 897 3533 920
rect 3571 939 3591 942
rect 3571 933 3574 939
rect 3588 933 3591 939
rect 3552 912 3555 915
rect 3552 909 3570 912
rect 3580 902 3583 909
rect 3580 899 3597 902
rect 3502 896 3521 897
rect 3497 894 3521 896
rect 3530 894 3573 897
rect 3503 888 3506 894
rect 3594 888 3597 899
rect 3559 883 3584 886
rect 3594 884 3607 888
rect 3559 881 3562 883
rect 3473 865 3489 868
rect 3494 865 3504 868
rect 3512 868 3515 876
rect 3524 878 3562 881
rect 3594 880 3597 884
rect 3524 868 3527 878
rect 3565 877 3597 880
rect 3565 874 3568 877
rect 3512 865 3527 868
rect 3512 862 3515 865
rect 3564 871 3570 874
rect 3503 852 3506 856
rect 3524 855 3529 858
rect 3542 858 3545 862
rect 3589 858 3592 862
rect 3534 855 3598 858
rect 3524 852 3527 855
rect 3497 849 3527 852
rect 3603 851 3607 884
rect 3603 844 3607 846
rect 3505 805 3533 808
rect 3506 799 3509 805
rect 3530 804 3533 805
rect 3530 801 3601 804
rect 3473 775 3492 778
rect 3497 776 3507 779
rect 3515 779 3518 787
rect 3545 795 3548 801
rect 3564 795 3567 801
rect 3515 776 3536 779
rect 3515 773 3518 776
rect 3506 763 3509 767
rect 3500 761 3524 763
rect 3500 760 3518 761
rect 3523 760 3524 761
rect 3533 753 3536 776
rect 3574 795 3594 798
rect 3574 789 3577 795
rect 3591 789 3594 795
rect 3555 768 3558 771
rect 3555 765 3573 768
rect 3583 758 3586 765
rect 3583 755 3600 758
rect 3505 752 3524 753
rect 3500 750 3524 752
rect 3533 750 3576 753
rect 3506 744 3509 750
rect 3597 744 3600 755
rect 3562 739 3587 742
rect 3597 740 3610 744
rect 3562 737 3565 739
rect 3473 721 3492 724
rect 3497 721 3507 724
rect 3515 724 3518 732
rect 3527 734 3565 737
rect 3597 736 3600 740
rect 3527 724 3530 734
rect 3568 733 3600 736
rect 3568 730 3571 733
rect 3515 721 3530 724
rect 3515 718 3518 721
rect 3567 727 3573 730
rect 3506 708 3509 712
rect 3527 711 3532 714
rect 3545 714 3548 718
rect 3592 714 3595 718
rect 3537 711 3601 714
rect 3527 708 3530 711
rect 3500 705 3530 708
rect 3606 705 3610 740
rect 3512 680 3540 683
rect 3513 674 3516 680
rect 3537 679 3540 680
rect 3537 676 3608 679
rect 3473 650 3499 653
rect 3504 651 3514 654
rect 3522 654 3525 662
rect 3552 670 3555 676
rect 3571 670 3574 676
rect 3522 651 3543 654
rect 3522 648 3525 651
rect 3513 638 3516 642
rect 3507 636 3531 638
rect 3507 635 3525 636
rect 3530 635 3531 636
rect 3540 628 3543 651
rect 3581 670 3601 673
rect 3581 664 3584 670
rect 3598 664 3601 670
rect 3562 643 3565 646
rect 3562 640 3580 643
rect 3590 633 3593 640
rect 3590 630 3607 633
rect 3512 627 3531 628
rect 3507 625 3531 627
rect 3540 625 3583 628
rect 3513 619 3516 625
rect 3604 619 3607 630
rect 3569 614 3594 617
rect 3604 615 3617 619
rect 3569 612 3572 614
rect 3473 596 3499 599
rect 3504 596 3514 599
rect 3522 599 3525 607
rect 3534 609 3572 612
rect 3604 611 3607 615
rect 3534 599 3537 609
rect 3575 608 3607 611
rect 3575 605 3578 608
rect 3522 596 3537 599
rect 3522 593 3525 596
rect 3574 602 3580 605
rect 3513 583 3516 587
rect 3534 586 3539 589
rect 3552 589 3555 593
rect 3599 589 3602 593
rect 3544 586 3608 589
rect 3534 583 3537 586
rect 3507 580 3537 583
rect 3613 578 3617 615
rect 3535 460 3558 464
rect 3539 458 3558 460
rect 3535 449 3539 454
rect 3554 449 3558 458
rect 3571 453 3595 454
rect 3571 449 3587 453
rect 3591 449 3595 453
rect 3571 447 3595 449
rect 3577 442 3581 447
rect 3546 421 3550 429
rect 3546 417 3558 421
rect 3554 415 3558 417
rect 3585 415 3589 422
rect 3473 410 3547 414
rect 3554 411 3578 415
rect 3585 411 3608 415
rect 3473 403 3536 407
rect 3554 400 3558 411
rect 3585 408 3589 411
rect 3592 410 3608 411
rect 3577 394 3581 398
rect 3571 393 3596 394
rect 3571 389 3591 393
rect 3571 388 3596 389
rect 3535 376 3539 380
rect 3535 372 3551 376
rect 3706 372 3709 1446
rect 3858 1447 3868 1450
rect 3876 1450 3879 1458
rect 3906 1466 3909 1472
rect 3925 1466 3928 1472
rect 3876 1447 3897 1450
rect 3876 1444 3879 1447
rect 3867 1434 3870 1438
rect 3861 1432 3885 1434
rect 3861 1431 3879 1432
rect 3884 1431 3885 1432
rect 3894 1424 3897 1447
rect 3935 1466 3955 1469
rect 3935 1460 3938 1466
rect 3952 1460 3955 1466
rect 3916 1439 3919 1442
rect 3916 1436 3934 1439
rect 3944 1429 3947 1436
rect 3944 1426 3961 1429
rect 3866 1423 3885 1424
rect 3861 1421 3885 1423
rect 3894 1421 3937 1424
rect 3867 1415 3870 1421
rect 3958 1415 3961 1426
rect 3923 1410 3948 1413
rect 3958 1411 3971 1415
rect 3923 1408 3926 1410
rect 3785 1392 3853 1397
rect 3858 1392 3868 1395
rect 3876 1395 3879 1403
rect 3888 1405 3926 1408
rect 3958 1407 3961 1411
rect 3888 1395 3891 1405
rect 3929 1404 3961 1407
rect 3967 1404 3971 1411
rect 3929 1401 3932 1404
rect 3876 1392 3891 1395
rect 3876 1389 3879 1392
rect 3928 1398 3934 1401
rect 3967 1400 3976 1404
rect 3867 1379 3870 1383
rect 3888 1382 3893 1385
rect 3906 1385 3909 1389
rect 3953 1385 3956 1389
rect 3898 1382 3962 1385
rect 3888 1379 3891 1382
rect 3861 1376 3891 1379
rect 3961 1296 3984 1300
rect 3961 1219 3965 1296
rect 3929 1215 3965 1219
rect 3869 1176 3872 1210
rect 3929 1209 3933 1215
rect 3915 1206 3940 1209
rect 3875 1200 3884 1203
rect 3875 1186 3878 1200
rect 3915 1195 3918 1206
rect 3908 1192 3918 1195
rect 3875 1183 3884 1186
rect 3869 1173 3878 1176
rect 3869 1157 3872 1173
rect 3905 1167 3908 1182
rect 3902 1164 3908 1167
rect 3869 1154 3878 1157
rect 3869 1142 3872 1154
rect 3920 1145 3923 1185
rect 3931 1174 3934 1196
rect 3937 1180 3940 1206
rect 3959 1204 3962 1210
rect 3955 1201 3962 1204
rect 3943 1180 3946 1182
rect 3937 1177 3946 1180
rect 3943 1176 3946 1177
rect 3931 1171 3939 1174
rect 3865 1139 3872 1142
rect 3894 1142 3923 1145
rect 3865 1118 3868 1139
rect 3894 1127 3897 1142
rect 3936 1139 3939 1171
rect 3959 1157 3962 1201
rect 4098 1167 4148 1171
rect 3955 1154 3962 1157
rect 3959 1146 3962 1154
rect 3959 1139 3962 1141
rect 3936 1136 3952 1139
rect 3959 1136 3968 1139
rect 3910 1132 3913 1133
rect 3910 1127 3912 1132
rect 3886 1124 3900 1127
rect 3865 1115 3874 1118
rect 3865 1114 3868 1115
rect 3894 1106 3897 1116
rect 3910 1118 3913 1127
rect 3906 1115 3913 1118
rect 3910 1109 3913 1115
rect 3920 1118 3923 1133
rect 3949 1127 3952 1136
rect 3941 1124 3955 1127
rect 3920 1115 3929 1118
rect 3920 1114 3923 1115
rect 3921 1109 3923 1114
rect 3949 1106 3952 1116
rect 3965 1118 3968 1136
rect 3961 1115 3968 1118
rect 3965 1109 3968 1115
rect 4038 1128 4041 1162
rect 4098 1161 4102 1167
rect 4084 1158 4109 1161
rect 4044 1152 4053 1155
rect 4044 1138 4047 1152
rect 4084 1147 4087 1158
rect 4077 1144 4087 1147
rect 4044 1135 4053 1138
rect 4038 1125 4047 1128
rect 4038 1109 4041 1125
rect 4074 1119 4077 1134
rect 4071 1116 4077 1119
rect 4038 1106 4047 1109
rect 3830 897 3834 913
rect 3895 905 3898 1101
rect 3949 1078 3952 1101
rect 4038 1094 4041 1106
rect 4089 1097 4092 1137
rect 4100 1126 4103 1148
rect 4106 1132 4109 1158
rect 4128 1156 4131 1162
rect 4124 1153 4131 1156
rect 4112 1132 4115 1134
rect 4106 1129 4115 1132
rect 4112 1128 4115 1129
rect 4100 1123 4108 1126
rect 4034 1091 4041 1094
rect 4063 1094 4092 1097
rect 3948 1075 3953 1078
rect 4034 1070 4037 1091
rect 4063 1079 4066 1094
rect 4105 1091 4108 1123
rect 4128 1109 4131 1153
rect 4124 1106 4131 1109
rect 4128 1098 4131 1106
rect 4128 1091 4131 1093
rect 4105 1088 4121 1091
rect 4128 1088 4137 1091
rect 4079 1084 4082 1085
rect 4079 1079 4081 1084
rect 4055 1076 4069 1079
rect 4034 1067 4043 1070
rect 4034 1066 4037 1067
rect 4063 1058 4066 1068
rect 4079 1070 4082 1079
rect 4075 1067 4082 1070
rect 4079 1061 4082 1067
rect 4089 1070 4092 1085
rect 4118 1079 4121 1088
rect 4110 1076 4124 1079
rect 4089 1067 4098 1070
rect 4089 1066 4092 1067
rect 4090 1061 4092 1066
rect 4118 1058 4121 1068
rect 4134 1070 4137 1088
rect 4130 1067 4137 1070
rect 4134 1061 4137 1067
rect 3887 901 3905 905
rect 3830 893 3847 897
rect 3934 897 3938 913
rect 3925 893 3938 897
rect 3837 892 3841 893
rect 3837 887 3841 888
rect 3798 643 3803 644
rect 3798 638 3803 639
rect 3789 634 3809 638
rect 3798 620 3803 634
rect 3897 630 3901 861
rect 3997 854 4001 874
rect 4064 862 4067 1053
rect 4118 1048 4121 1053
rect 4281 1009 4326 1013
rect 4221 970 4224 1004
rect 4281 1003 4285 1009
rect 4267 1000 4292 1003
rect 4227 994 4236 997
rect 4227 980 4230 994
rect 4267 989 4270 1000
rect 4260 986 4270 989
rect 4227 977 4236 980
rect 4221 967 4230 970
rect 4221 951 4224 967
rect 4257 961 4260 976
rect 4254 958 4260 961
rect 4221 948 4230 951
rect 4221 936 4224 948
rect 4272 939 4275 979
rect 4283 968 4286 990
rect 4289 974 4292 1000
rect 4311 998 4314 1004
rect 4307 995 4314 998
rect 4295 974 4298 976
rect 4289 971 4298 974
rect 4295 970 4298 971
rect 4283 965 4291 968
rect 4217 933 4224 936
rect 4246 936 4275 939
rect 4217 912 4220 933
rect 4246 921 4249 936
rect 4288 933 4291 965
rect 4311 951 4314 995
rect 4307 948 4314 951
rect 4311 940 4314 948
rect 4311 933 4314 935
rect 4288 930 4304 933
rect 4311 930 4320 933
rect 4262 926 4265 927
rect 4262 921 4264 926
rect 4238 918 4252 921
rect 4217 909 4226 912
rect 4217 908 4220 909
rect 4246 900 4249 910
rect 4262 912 4265 921
rect 4258 909 4265 912
rect 4262 903 4265 909
rect 4272 912 4275 927
rect 4301 921 4304 930
rect 4293 918 4307 921
rect 4272 909 4281 912
rect 4272 908 4275 909
rect 4273 903 4275 908
rect 4301 900 4304 910
rect 4317 912 4320 930
rect 4313 909 4320 912
rect 4317 903 4320 909
rect 4054 858 4072 862
rect 3997 850 4014 854
rect 4101 854 4105 874
rect 4092 850 4105 854
rect 3997 843 4001 850
rect 4004 849 4008 850
rect 4004 844 4008 845
rect 4101 843 4105 850
rect 4179 847 4183 863
rect 4247 855 4250 895
rect 4301 892 4304 895
rect 4301 886 4306 892
rect 4236 851 4254 855
rect 4179 843 4196 847
rect 4283 847 4287 863
rect 4274 843 4287 847
rect 4179 835 4183 843
rect 4186 842 4190 843
rect 4186 837 4190 838
rect 4283 835 4287 843
rect 4064 811 4069 817
rect 3972 666 3977 667
rect 3972 661 3977 662
rect 3963 657 3983 661
rect 3972 643 3977 657
rect 4065 653 4069 811
rect 4246 800 4251 804
rect 4247 785 4250 800
rect 4146 670 4151 671
rect 4146 665 4151 666
rect 4137 661 4157 665
rect 4033 649 4069 653
rect 3859 626 3901 630
rect 3897 589 3901 626
rect 4065 599 4069 649
rect 4146 647 4151 661
rect 4246 657 4250 785
rect 4474 772 4495 776
rect 4482 769 4486 772
rect 4476 765 4477 769
rect 4481 765 4486 769
rect 4482 759 4486 765
rect 4342 705 4347 706
rect 4436 704 4482 709
rect 4490 708 4494 719
rect 4490 704 4504 708
rect 4342 700 4347 701
rect 4333 696 4353 700
rect 4342 682 4347 696
rect 4436 692 4440 704
rect 4490 701 4494 704
rect 4403 688 4440 692
rect 4207 653 4250 657
rect 4246 607 4250 653
rect 4436 615 4440 688
rect 4482 672 4486 681
rect 4474 668 4491 672
rect 4429 611 4440 615
rect 4241 603 4329 607
rect 4064 597 4141 599
rect 4060 595 4141 597
rect 4060 593 4068 595
rect 3892 585 3960 589
rect 3690 367 3709 372
rect 3739 577 3792 581
rect 3739 471 3743 577
rect 3897 475 3901 585
rect 4064 486 4068 593
rect 4245 496 4249 603
rect 4436 506 4440 611
rect 4431 502 4440 506
rect 4239 492 4249 496
rect 4324 494 4331 498
rect 4059 482 4068 486
rect 4133 484 4139 488
rect 3891 471 3901 475
rect 3953 474 3959 478
rect 3785 463 3791 467
rect 3535 351 3558 355
rect 3539 349 3558 351
rect 3535 340 3539 345
rect 3554 340 3558 349
rect 3690 348 3695 367
rect 3706 364 3709 367
rect 3747 369 3751 371
rect 3786 458 3790 463
rect 3953 458 3957 474
rect 4133 458 4137 484
rect 4324 458 4328 494
rect 3786 454 4328 458
rect 3786 369 3790 454
rect 3924 373 3930 377
rect 3747 365 3824 369
rect 3571 344 3595 345
rect 3571 340 3587 344
rect 3591 340 3595 344
rect 3690 343 3730 348
rect 3571 338 3595 340
rect 3577 333 3581 338
rect 3546 312 3550 320
rect 3546 308 3558 312
rect 3554 306 3558 308
rect 3585 306 3589 313
rect 3680 309 3684 325
rect 3725 317 3730 343
rect 3864 338 3868 347
rect 3921 344 3931 346
rect 3936 344 3939 346
rect 3921 342 3939 344
rect 3864 334 3881 338
rect 3968 338 3972 343
rect 3959 334 3972 338
rect 3864 324 3868 334
rect 3871 333 3875 334
rect 3871 328 3875 329
rect 3968 325 3972 334
rect 3715 313 3737 317
rect 3473 301 3547 305
rect 3554 302 3578 306
rect 3585 302 3621 306
rect 3680 305 3690 309
rect 3752 309 3756 317
rect 3473 294 3536 298
rect 3554 291 3558 302
rect 3585 299 3589 302
rect 3577 285 3581 289
rect 3571 284 3596 285
rect 3571 280 3591 284
rect 3571 279 3596 280
rect 3535 267 3539 271
rect 3535 263 3551 267
rect 3680 264 3684 305
rect 3724 285 3729 306
rect 3747 305 3756 309
rect 3690 282 3747 285
rect 3690 272 3715 282
rect 3730 273 3734 274
rect 3737 274 3747 282
rect 3680 260 3690 264
rect 3536 232 3559 236
rect 3540 230 3559 232
rect 3536 221 3540 226
rect 3555 221 3559 230
rect 3572 225 3596 226
rect 3572 221 3588 225
rect 3592 221 3596 225
rect 3572 219 3596 221
rect 3680 220 3684 260
rect 3752 258 3756 305
rect 3747 254 3756 258
rect 3729 250 3734 254
rect 3724 246 3734 250
rect 3724 241 3729 246
rect 3690 238 3747 241
rect 3690 228 3715 238
rect 3730 229 3734 230
rect 3737 230 3747 238
rect 3578 214 3582 219
rect 3680 216 3690 220
rect 3547 193 3551 201
rect 3547 189 3559 193
rect 3555 187 3559 189
rect 3586 187 3590 194
rect 3473 182 3548 186
rect 3555 183 3579 187
rect 3586 183 3633 187
rect 3473 175 3537 179
rect 3555 172 3559 183
rect 3586 180 3590 183
rect 3680 182 3684 216
rect 3752 214 3756 254
rect 3747 210 3756 214
rect 3722 202 3726 203
rect 3729 207 3734 210
rect 3729 202 3731 207
rect 3715 194 3747 198
rect 3680 178 3690 182
rect 3730 178 3734 187
rect 3737 186 3747 194
rect 3752 178 3756 210
rect 3680 172 3684 178
rect 3578 166 3582 170
rect 3722 167 3726 174
rect 3747 174 3756 178
rect 3752 173 3756 174
rect 3572 165 3597 166
rect 3572 161 3592 165
rect 3572 160 3597 161
rect 3536 148 3540 152
rect 3536 144 3552 148
rect 3540 124 3563 128
rect 3544 122 3563 124
rect 3540 113 3544 118
rect 3559 113 3563 122
rect 3576 117 3600 118
rect 3576 113 3592 117
rect 3596 113 3600 117
rect 3576 111 3600 113
rect 3582 106 3586 111
rect 3551 85 3555 93
rect 3551 81 3563 85
rect 3559 79 3563 81
rect 3590 79 3594 86
rect 3473 74 3552 78
rect 3559 75 3583 79
rect 3590 75 3647 79
rect 3473 67 3541 71
rect 3559 64 3563 75
rect 3590 72 3594 75
rect 3582 58 3586 62
rect 3576 57 3601 58
rect 3576 53 3596 57
rect 3576 52 3601 53
rect 3540 40 3544 44
rect 3540 36 3556 40
<< m2contact >>
rect 3488 1050 3493 1055
rect 3488 996 3493 1001
rect 3602 976 3607 981
rect 3489 918 3494 923
rect 3489 864 3494 869
rect 3602 846 3607 851
rect 3492 774 3497 779
rect 3492 720 3497 725
rect 3606 700 3611 705
rect 3499 649 3504 654
rect 3499 595 3504 600
rect 3613 573 3618 578
rect 3608 410 3613 415
rect 3853 1445 3858 1450
rect 3780 1392 3785 1397
rect 3853 1391 3858 1396
rect 3894 1101 3899 1106
rect 3948 1101 3953 1106
rect 3948 1070 3953 1075
rect 4063 1053 4068 1058
rect 4117 1053 4122 1058
rect 3897 861 3902 867
rect 4118 1042 4124 1048
rect 4246 895 4251 900
rect 4300 895 4305 900
rect 4301 880 4306 886
rect 4064 817 4069 825
rect 4246 804 4251 810
rect 3706 359 3711 364
rect 3931 344 3936 349
rect 3621 302 3626 307
rect 3729 274 3734 279
rect 3729 230 3734 235
rect 3633 183 3639 189
rect 3721 203 3726 208
rect 3731 202 3736 207
rect 3729 173 3734 178
rect 3647 75 3652 81
<< pm12contact >>
rect 3544 1033 3549 1038
rect 3553 1032 3558 1037
rect 3545 901 3550 906
rect 3554 900 3559 905
rect 3548 757 3553 762
rect 3557 756 3562 761
rect 3555 632 3560 637
rect 3564 631 3569 636
rect 3909 1428 3914 1433
rect 3918 1427 3923 1432
rect 3912 1166 3917 1171
rect 3911 1157 3916 1162
rect 4081 1118 4086 1123
rect 4080 1109 4085 1114
rect 3897 893 3902 898
rect 3876 633 3882 639
rect 4264 960 4269 965
rect 4263 951 4268 956
rect 4064 850 4069 855
rect 4246 843 4251 848
rect 4050 656 4056 662
rect 4224 660 4230 666
rect 4420 695 4426 701
rect 4317 610 4322 615
rect 4129 602 4134 607
rect 3948 592 3953 597
rect 3780 584 3785 589
rect 4319 501 4324 506
rect 4127 491 4132 496
rect 3947 481 3952 486
rect 3779 470 3784 475
rect 3931 365 3936 370
rect 3739 359 3744 364
rect 3931 334 3936 339
<< metal2 >>
rect 3854 1439 3857 1445
rect 3854 1436 3891 1439
rect 3888 1433 3891 1436
rect 3888 1430 3909 1433
rect 3918 1417 3921 1427
rect 3855 1414 3921 1417
rect 3855 1396 3858 1414
rect 3489 1044 3492 1050
rect 3489 1041 3526 1044
rect 3523 1038 3526 1041
rect 3523 1035 3544 1038
rect 3553 1022 3556 1032
rect 3490 1019 3556 1022
rect 3490 1001 3493 1019
rect 3607 976 3662 981
rect 3490 912 3493 918
rect 3490 909 3527 912
rect 3524 906 3527 909
rect 3524 903 3545 906
rect 3554 890 3557 900
rect 3491 887 3557 890
rect 3491 869 3494 887
rect 3607 846 3650 851
rect 3493 768 3496 774
rect 3493 765 3530 768
rect 3527 762 3530 765
rect 3527 759 3548 762
rect 3557 746 3560 756
rect 3494 743 3560 746
rect 3494 725 3497 743
rect 3611 701 3629 705
rect 3500 643 3503 649
rect 3500 640 3537 643
rect 3534 637 3537 640
rect 3534 634 3555 637
rect 3564 621 3567 631
rect 3501 618 3567 621
rect 3501 600 3504 618
rect 3613 537 3618 573
rect 3625 547 3629 701
rect 3645 557 3650 846
rect 3657 572 3662 976
rect 3780 597 3785 1392
rect 3917 1166 3930 1169
rect 3911 1139 3914 1157
rect 3905 1136 3914 1139
rect 3905 1105 3908 1136
rect 3899 1102 3908 1105
rect 3927 1106 3930 1166
rect 4086 1118 4099 1121
rect 3927 1103 3948 1106
rect 4080 1091 4083 1109
rect 4074 1088 4083 1091
rect 3897 867 3902 893
rect 3876 639 3882 643
rect 3948 607 3953 1070
rect 4074 1057 4077 1088
rect 4068 1054 4077 1057
rect 4096 1058 4099 1118
rect 4096 1055 4117 1058
rect 4124 1042 4133 1046
rect 4064 825 4069 850
rect 4050 662 4056 666
rect 4129 616 4133 1042
rect 4269 960 4282 963
rect 4263 933 4266 951
rect 4257 930 4266 933
rect 4257 899 4260 930
rect 4251 896 4260 899
rect 4279 900 4282 960
rect 4279 897 4300 900
rect 4246 810 4251 843
rect 4301 791 4306 880
rect 4301 786 4322 791
rect 4301 785 4306 786
rect 4224 666 4230 670
rect 4317 628 4322 786
rect 4420 701 4426 705
rect 3770 592 3785 597
rect 3770 572 3775 592
rect 3780 589 3785 592
rect 3939 602 3953 607
rect 3657 567 3775 572
rect 3939 557 3944 602
rect 3948 597 3953 602
rect 4120 612 4133 616
rect 3645 552 3944 557
rect 4120 547 4124 612
rect 4129 611 4133 612
rect 4304 623 4322 628
rect 4129 607 4134 611
rect 3625 543 4124 547
rect 4304 537 4309 623
rect 4317 615 4322 623
rect 3613 532 4309 537
rect 3608 508 4324 513
rect 3608 415 3613 508
rect 4319 506 4324 508
rect 3621 498 4132 503
rect 3621 307 3626 498
rect 4127 496 4132 498
rect 3633 487 3952 493
rect 3633 189 3639 487
rect 3947 486 3952 487
rect 3647 478 3784 483
rect 3647 81 3652 478
rect 3779 475 3784 478
rect 3711 359 3739 364
rect 3931 359 3936 365
rect 3931 349 3936 354
rect 3931 331 3936 334
rect 3758 279 3761 283
rect 3734 274 3761 279
rect 3673 230 3729 234
rect 3673 207 3677 230
rect 3673 203 3721 207
rect 3758 207 3761 274
rect 3736 203 3761 207
rect 3730 170 3734 173
rect 3758 170 3761 203
rect 3730 164 3761 170
rect 3730 152 3734 164
<< m3contact >>
rect 3876 643 3882 649
rect 4050 666 4056 672
rect 4224 670 4230 676
rect 4420 705 4426 711
rect 3931 354 3936 359
<< m123contact >>
rect 3861 1476 3866 1481
rect 3861 1423 3866 1428
rect 3879 1427 3884 1432
rect 3496 1081 3501 1086
rect 3496 1028 3501 1033
rect 3514 1032 3519 1037
rect 3528 987 3533 992
rect 3497 949 3502 954
rect 3497 896 3502 901
rect 3515 900 3520 905
rect 3529 855 3534 860
rect 3500 805 3505 810
rect 3500 752 3505 757
rect 3518 756 3523 761
rect 3532 711 3537 716
rect 3507 680 3512 685
rect 3507 627 3512 632
rect 3525 631 3530 636
rect 3539 586 3544 591
rect 3893 1382 3898 1387
rect 3863 1109 3868 1114
rect 3912 1127 3917 1132
rect 3916 1109 3921 1114
rect 3957 1141 3962 1146
rect 4032 1061 4037 1066
rect 4081 1079 4086 1084
rect 4085 1061 4090 1066
rect 4126 1093 4131 1098
rect 4215 903 4220 908
rect 4264 921 4269 926
rect 4268 903 4273 908
rect 4309 935 4314 940
<< metal3 >>
rect 3861 1428 3864 1476
rect 3884 1427 3896 1430
rect 3893 1387 3896 1427
rect 3914 1141 3957 1144
rect 3914 1132 3917 1141
rect 3868 1109 3916 1112
rect 4083 1093 4126 1096
rect 4083 1084 4086 1093
rect 3496 1033 3499 1081
rect 4037 1061 4085 1064
rect 3519 1032 3531 1035
rect 3528 992 3531 1032
rect 3497 901 3500 949
rect 4266 935 4309 938
rect 4266 926 4269 935
rect 4220 903 4268 906
rect 3520 900 3532 903
rect 3529 860 3532 900
rect 3500 757 3503 805
rect 3523 756 3535 759
rect 3532 716 3535 756
rect 3876 736 4426 741
rect 3507 632 3510 680
rect 3876 649 3882 736
rect 4050 672 4056 736
rect 3530 631 3542 634
rect 3539 591 3542 631
rect 4088 359 4093 736
rect 4224 676 4230 736
rect 4420 711 4426 736
rect 3936 354 4093 359
<< labels >>
rlabel metal1 3894 471 3899 475 3 pdr1
rlabel metal2 3779 475 3784 479 3 gen_1
rlabel metal1 3739 474 3743 479 1 prop1_car0
rlabel metal2 3735 359 3739 364 1 carry_0
rlabel metal1 3747 365 3751 370 1 clock_car0
rlabel metal1 3816 365 3821 369 7 clock_car0
rlabel metal2 3931 361 3936 365 7 clock_in
rlabel metal1 3925 373 3930 377 7 gnd!
rlabel metal1 3785 463 3790 467 3 clock_car0
rlabel metal1 3896 585 3900 589 3 pdr1
rlabel metal2 3780 589 3785 593 4 prop_1
rlabel metal1 3786 577 3791 581 3 prop1_car0
rlabel metal1 3789 634 3794 638 3 vdd!
rlabel m3contact 3876 643 3882 649 6 clock_in
rlabel metal1 3868 626 3873 630 7 pdr1
rlabel metal1 3953 474 3958 478 3 clock_car0
rlabel metal2 3947 486 3952 490 3 gen_2
rlabel metal1 4062 482 4067 486 3 pdr2
rlabel metal1 4063 593 4068 597 3 pdr2
rlabel metal2 3948 597 3953 601 3 prop_2
rlabel metal1 3954 585 3959 589 3 pdr1
rlabel metal1 3963 657 3968 661 3 vdd!
rlabel m3contact 4050 666 4056 672 7 clock_in
rlabel metal1 4043 649 4047 653 7 pdr2
rlabel metal1 4133 484 4138 488 3 clock_car0
rlabel metal2 4127 496 4132 500 3 gen_3
rlabel metal1 4242 492 4247 496 3 pdr3
rlabel metal1 4434 502 4439 506 3 pdr4
rlabel metal2 4319 506 4324 510 3 gen_4
rlabel metal1 4325 494 4330 498 1 clock_car0
rlabel metal1 4244 603 4249 607 3 pdr3
rlabel metal2 4129 607 4134 611 3 prop_3
rlabel metal1 4135 595 4140 599 3 pdr2
rlabel metal1 4432 611 4437 615 3 pdr4
rlabel metal2 4317 615 4322 619 3 prop_4
rlabel metal1 4323 603 4328 607 3 pdr3
rlabel metal1 4137 661 4142 665 3 vdd!
rlabel m3contact 4224 670 4230 676 7 clock_in
rlabel metal1 4217 653 4221 657 7 pdr3
rlabel metal1 4333 696 4338 700 3 vdd!
rlabel m3contact 4420 706 4426 711 7 clock_in
rlabel metal1 4413 688 4417 692 7 pdr4
rlabel metal1 4490 704 4494 709 1 c4
rlabel metal1 4483 772 4488 776 5 vdd!
rlabel metal1 4487 668 4491 672 1 gnd!
rlabel metal1 3968 339 3972 343 7 gnd!
rlabel metal1 3864 335 3868 340 3 vdd!
rlabel metal2 3931 331 3936 334 7 clk_org
rlabel metal1 3931 342 3936 346 7 clock_in
rlabel metal1 3970 1413 3970 1413 1 s1
rlabel metal1 3851 1394 3851 1394 1 prop_1
rlabel metal1 3851 1448 3851 1448 1 carry_0
rlabel metal1 3874 1422 3877 1424 1 vdd
rlabel metal1 3873 1476 3876 1478 5 vdd
rlabel metal1 3877 1432 3878 1434 1 gnd
rlabel metal1 3929 1382 3932 1384 1 gnd
rlabel metal1 3879 1376 3883 1379 1 gnd
rlabel metal1 3550 125 3550 125 5 vdd
rlabel metal1 3551 38 3551 38 1 gnd
rlabel metal1 3583 56 3583 56 1 gnd
rlabel metal1 3580 113 3580 113 5 vdd
rlabel metal1 3535 76 3535 76 3 q_a1
rlabel metal1 3537 69 3537 69 3 q_b1
rlabel metal1 3599 76 3599 76 1 gen_1
rlabel metal1 3546 233 3546 233 5 vdd
rlabel metal1 3547 146 3547 146 1 gnd
rlabel metal1 3579 164 3579 164 1 gnd
rlabel metal1 3576 221 3576 221 5 vdd
rlabel metal1 3532 183 3532 183 1 q_a2
rlabel metal1 3532 176 3532 176 1 q_b2
rlabel metal1 3595 185 3595 185 1 gen_2
rlabel metal1 3545 352 3545 352 5 vdd
rlabel metal1 3546 265 3546 265 1 gnd
rlabel metal1 3578 283 3578 283 1 gnd
rlabel metal1 3575 340 3575 340 5 vdd
rlabel metal1 3530 302 3530 302 1 q_b3
rlabel metal1 3532 295 3532 295 1 q_a3
rlabel metal1 3593 304 3593 304 1 gen_3
rlabel metal1 3545 461 3545 461 5 vdd
rlabel metal1 3546 374 3546 374 1 gnd
rlabel metal1 3578 392 3578 392 1 gnd
rlabel metal1 3575 449 3575 449 5 vdd
rlabel metal1 3530 412 3530 412 3 q_a4
rlabel metal1 3530 406 3530 406 3 q_b4
rlabel metal1 3593 413 3593 413 1 gen_4
rlabel metal1 3605 887 3605 887 1 prop_2
rlabel metal1 3487 866 3487 866 3 q_b2
rlabel metal1 3487 921 3487 921 3 q_a2
rlabel metal1 3510 895 3513 897 1 vdd
rlabel metal1 3509 949 3512 951 5 vdd
rlabel metal1 3513 905 3514 907 1 gnd
rlabel metal1 3565 855 3568 857 1 gnd
rlabel metal1 3515 849 3519 852 1 gnd
rlabel metal1 3518 705 3522 708 1 gnd
rlabel metal1 3568 711 3571 713 1 gnd
rlabel metal1 3516 761 3517 763 1 gnd
rlabel metal1 3512 805 3515 807 5 vdd
rlabel metal1 3513 751 3516 753 1 vdd
rlabel metal1 3491 777 3491 777 1 q_a3
rlabel metal1 3491 723 3491 723 1 q_b3
rlabel metal1 3608 742 3608 742 1 prop_3
rlabel metal1 3525 580 3529 583 1 gnd
rlabel metal1 3575 586 3578 588 1 gnd
rlabel metal1 3523 636 3524 638 1 gnd
rlabel metal1 3519 680 3522 682 5 vdd
rlabel metal1 3520 626 3523 628 1 vdd
rlabel metal1 3497 651 3497 651 1 q_a4
rlabel metal1 3497 598 3497 598 1 q_b4
rlabel metal1 3616 617 3616 617 1 prop_4
rlabel metal1 3602 1018 3602 1018 1 prop_1
rlabel metal1 3486 999 3486 999 1 q_b1
rlabel metal1 3486 1053 3486 1053 1 q_a1
rlabel metal1 3509 1027 3512 1029 1 vdd
rlabel metal1 3508 1081 3511 1083 5 vdd
rlabel metal1 3512 1037 3513 1039 1 gnd
rlabel metal1 3564 987 3567 989 1 gnd
rlabel metal1 3514 981 3518 984 1 gnd
rlabel metal1 3753 182 3754 185 7 gnd
rlabel metal1 3681 188 3682 190 3 vdd
rlabel metal2 3733 169 3733 169 7 clk_org
rlabel metal1 3724 168 3724 168 7 cin
rlabel metal1 3728 325 3728 325 7 carry_0
rlabel metal1 4249 893 4249 893 7 c3
rlabel metal1 4302 893 4302 893 7 prop_4
rlabel metal1 4283 1011 4283 1011 7 s4
rlabel metal1 4272 916 4274 919 7 vdd
rlabel metal1 4218 915 4220 918 3 vdd
rlabel metal1 4262 919 4264 920 7 gnd
rlabel metal1 4312 971 4314 974 7 gnd
rlabel metal1 4317 921 4320 925 7 gnd
rlabel metal2 4246 840 4251 843 7 pdr3
rlabel metal1 4246 851 4251 855 7 c3
rlabel metal1 4179 843 4183 847 3 vdd!
rlabel metal1 4283 847 4287 851 7 gnd!
rlabel metal1 3965 1127 3968 1131 7 gnd
rlabel metal1 3960 1177 3962 1180 7 gnd
rlabel metal1 3910 1125 3912 1126 7 gnd
rlabel metal1 3866 1121 3868 1124 3 vdd
rlabel metal1 3920 1122 3922 1125 7 vdd
rlabel metal1 3897 1100 3897 1100 7 c1
rlabel metal1 3951 1099 3951 1099 7 prop_2
rlabel metal1 3932 1218 3932 1218 5 s2
rlabel metal1 4134 1079 4137 1083 7 gnd
rlabel metal1 4129 1129 4131 1132 7 gnd
rlabel metal1 4079 1077 4081 1078 7 gnd
rlabel metal1 4035 1073 4037 1076 3 vdd
rlabel metal1 4089 1074 4091 1077 7 vdd
rlabel metal1 4065 1051 4065 1051 7 c2
rlabel metal1 4100 1170 4100 1170 7 s3
rlabel metal1 4120 1049 4120 1049 7 prop_3
rlabel metal1 3934 902 3938 906 7 gnd!
rlabel metal1 3830 893 3834 897 3 vdd!
rlabel metal1 3897 901 3902 905 7 c1
rlabel metal2 3897 890 3902 893 7 pdr1
rlabel metal1 4101 861 4105 865 7 gnd!
rlabel metal1 3997 850 4001 854 3 vdd!
rlabel metal1 4064 858 4069 862 7 c2
rlabel metal2 4064 847 4069 850 7 pdr2
<< end >>
