magic
tech scmos
timestamp 1732016630
<< nwell >>
rect 7996 2430 8028 2467
rect 8034 2430 8060 2467
rect 8078 2430 8104 2467
rect 8123 2430 8149 2467
rect 7990 2261 8022 2298
rect 8028 2261 8054 2298
rect 8072 2261 8098 2298
rect 8117 2261 8143 2298
rect 12487 2221 12511 2245
rect 12526 2235 12560 2241
rect 12526 2205 12588 2235
rect 12554 2199 12588 2205
rect 12487 2166 12511 2190
rect 7990 2081 8022 2118
rect 8028 2081 8054 2118
rect 8072 2081 8098 2118
rect 8117 2081 8143 2118
rect 8525 2084 8549 2108
rect 8564 2098 8598 2104
rect 8564 2068 8626 2098
rect 8592 2062 8626 2068
rect 8525 2029 8549 2053
rect 13402 2027 13426 2059
rect 10223 1948 10247 2010
rect 10273 1949 10297 2011
rect 10323 1949 10347 2011
rect 10370 1949 10394 2011
rect 12917 1967 12949 2004
rect 12955 1967 12981 2004
rect 12999 1967 13025 2004
rect 13044 1967 13070 2004
rect 9012 1870 9048 1910
rect 9054 1863 9078 1903
rect 8038 1765 8070 1802
rect 8076 1765 8102 1802
rect 8120 1765 8146 1802
rect 8165 1765 8191 1802
rect 8516 1725 8540 1749
rect 8555 1739 8589 1745
rect 8555 1709 8617 1739
rect 10692 1727 10716 1779
rect 10730 1727 10754 1779
rect 10774 1727 10798 1779
rect 10812 1727 10836 1779
rect 10858 1729 10882 1781
rect 8583 1703 8617 1709
rect 8516 1670 8540 1694
rect 8042 1603 8074 1640
rect 8080 1603 8106 1640
rect 8124 1603 8150 1640
rect 8169 1603 8195 1640
rect 13430 1606 13454 1638
rect 9014 1520 9050 1560
rect 9056 1513 9080 1553
rect 12902 1526 12934 1563
rect 12940 1526 12966 1563
rect 12984 1526 13010 1563
rect 13029 1526 13055 1563
rect 12527 1411 12551 1435
rect 12566 1425 12600 1431
rect 12566 1395 12628 1425
rect 8047 1353 8079 1390
rect 8085 1353 8111 1390
rect 8129 1353 8155 1390
rect 8174 1353 8200 1390
rect 8543 1366 8567 1390
rect 12594 1389 12628 1395
rect 8582 1380 8616 1386
rect 8582 1350 8644 1380
rect 12527 1356 12551 1380
rect 8610 1344 8644 1350
rect 8543 1311 8567 1335
rect 8045 1193 8077 1230
rect 8083 1193 8109 1230
rect 8127 1193 8153 1230
rect 8172 1193 8198 1230
rect 9022 1228 9058 1268
rect 9064 1221 9088 1261
rect 13481 1052 13505 1084
rect 8536 1023 8560 1047
rect 8575 1037 8609 1043
rect 8575 1007 8637 1037
rect 8603 1001 8637 1007
rect 8073 958 8105 995
rect 8111 958 8137 995
rect 8155 958 8181 995
rect 8200 958 8226 995
rect 8536 968 8560 992
rect 12467 981 12491 1005
rect 12506 995 12540 1001
rect 12506 965 12568 995
rect 12887 973 12919 1010
rect 12925 973 12951 1010
rect 12969 973 12995 1010
rect 13014 973 13040 1010
rect 12534 959 12568 965
rect 12467 926 12491 950
rect 8082 833 8114 870
rect 8120 833 8146 870
rect 8164 833 8190 870
rect 8209 833 8235 870
rect 9010 862 9046 902
rect 9052 855 9076 895
rect 12900 681 12932 718
rect 12938 681 12964 718
rect 12982 681 13008 718
rect 13027 681 13053 718
rect 13466 703 13490 735
rect 12424 445 12448 469
rect 12463 459 12497 465
rect 12463 429 12525 459
rect 12491 423 12525 429
rect 12424 390 12448 414
rect 12922 307 12954 344
rect 12960 307 12986 344
rect 13004 307 13030 344
rect 13049 307 13075 344
rect 13519 318 13543 350
<< ntransistor >>
rect 8003 2404 8005 2414
rect 8039 2404 8041 2414
rect 8047 2404 8049 2414
rect 8083 2404 8085 2414
rect 8091 2404 8093 2414
rect 8134 2404 8136 2414
rect 7997 2235 7999 2245
rect 8033 2235 8035 2245
rect 8041 2235 8043 2245
rect 8077 2235 8079 2245
rect 8085 2235 8087 2245
rect 8128 2235 8130 2245
rect 12498 2207 12500 2213
rect 12537 2158 12539 2170
rect 12547 2158 12549 2170
rect 12565 2158 12567 2170
rect 12575 2158 12577 2170
rect 12498 2152 12500 2158
rect 8536 2070 8538 2076
rect 7997 2055 7999 2065
rect 8033 2055 8035 2065
rect 8041 2055 8043 2065
rect 8077 2055 8079 2065
rect 8085 2055 8087 2065
rect 8128 2055 8130 2065
rect 8575 2021 8577 2033
rect 8585 2021 8587 2033
rect 8603 2021 8605 2033
rect 8613 2021 8615 2033
rect 8536 2015 8538 2021
rect 13413 2005 13415 2015
rect 12924 1941 12926 1951
rect 12960 1941 12962 1951
rect 12968 1941 12970 1951
rect 13004 1941 13006 1951
rect 13012 1941 13014 1951
rect 13055 1941 13057 1951
rect 9023 1827 9025 1847
rect 9034 1827 9036 1847
rect 9065 1845 9067 1855
rect 8045 1739 8047 1749
rect 8081 1739 8083 1749
rect 8089 1739 8091 1749
rect 8125 1739 8127 1749
rect 8133 1739 8135 1749
rect 8176 1739 8178 1749
rect 8527 1711 8529 1717
rect 8566 1662 8568 1674
rect 8576 1662 8578 1674
rect 8594 1662 8596 1674
rect 8604 1662 8606 1674
rect 10170 1668 10172 1768
rect 10198 1668 10200 1768
rect 10225 1668 10227 1768
rect 10264 1668 10266 1768
rect 10292 1668 10294 1768
rect 10319 1668 10321 1768
rect 10359 1669 10361 1769
rect 10387 1669 10389 1769
rect 10414 1669 10416 1769
rect 10450 1669 10452 1769
rect 10703 1695 10705 1715
rect 10741 1695 10743 1715
rect 10785 1695 10787 1715
rect 10823 1695 10825 1715
rect 10869 1697 10871 1717
rect 8527 1656 8529 1662
rect 8049 1577 8051 1587
rect 8085 1577 8087 1587
rect 8093 1577 8095 1587
rect 8129 1577 8131 1587
rect 8137 1577 8139 1587
rect 8180 1577 8182 1587
rect 13441 1584 13443 1594
rect 9025 1477 9027 1497
rect 9036 1477 9038 1497
rect 9067 1495 9069 1505
rect 12909 1500 12911 1510
rect 12945 1500 12947 1510
rect 12953 1500 12955 1510
rect 12989 1500 12991 1510
rect 12997 1500 12999 1510
rect 13040 1500 13042 1510
rect 12538 1397 12540 1403
rect 8554 1352 8556 1358
rect 8054 1327 8056 1337
rect 8090 1327 8092 1337
rect 8098 1327 8100 1337
rect 8134 1327 8136 1337
rect 8142 1327 8144 1337
rect 8185 1327 8187 1337
rect 12577 1348 12579 1360
rect 12587 1348 12589 1360
rect 12605 1348 12607 1360
rect 12615 1348 12617 1360
rect 12538 1342 12540 1348
rect 8593 1303 8595 1315
rect 8603 1303 8605 1315
rect 8621 1303 8623 1315
rect 8631 1303 8633 1315
rect 8554 1297 8556 1303
rect 9033 1185 9035 1205
rect 9044 1185 9046 1205
rect 9075 1203 9077 1213
rect 8052 1167 8054 1177
rect 8088 1167 8090 1177
rect 8096 1167 8098 1177
rect 8132 1167 8134 1177
rect 8140 1167 8142 1177
rect 8183 1167 8185 1177
rect 8547 1009 8549 1015
rect 13492 1030 13494 1040
rect 8586 960 8588 972
rect 8596 960 8598 972
rect 8614 960 8616 972
rect 8624 960 8626 972
rect 12478 967 12480 973
rect 8547 954 8549 960
rect 8080 932 8082 942
rect 8116 932 8118 942
rect 8124 932 8126 942
rect 8160 932 8162 942
rect 8168 932 8170 942
rect 8211 932 8213 942
rect 12894 947 12896 957
rect 12930 947 12932 957
rect 12938 947 12940 957
rect 12974 947 12976 957
rect 12982 947 12984 957
rect 13025 947 13027 957
rect 12517 918 12519 930
rect 12527 918 12529 930
rect 12545 918 12547 930
rect 12555 918 12557 930
rect 12478 912 12480 918
rect 9021 819 9023 839
rect 9032 819 9034 839
rect 9063 837 9065 847
rect 8089 807 8091 817
rect 8125 807 8127 817
rect 8133 807 8135 817
rect 8169 807 8171 817
rect 8177 807 8179 817
rect 8220 807 8222 817
rect 13477 681 13479 691
rect 12907 655 12909 665
rect 12943 655 12945 665
rect 12951 655 12953 665
rect 12987 655 12989 665
rect 12995 655 12997 665
rect 13038 655 13040 665
rect 12435 431 12437 437
rect 12474 382 12476 394
rect 12484 382 12486 394
rect 12502 382 12504 394
rect 12512 382 12514 394
rect 12435 376 12437 382
rect 13530 296 13532 306
rect 12929 281 12931 291
rect 12965 281 12967 291
rect 12973 281 12975 291
rect 13009 281 13011 291
rect 13017 281 13019 291
rect 13060 281 13062 291
<< ptransistor >>
rect 8007 2436 8009 2461
rect 8015 2436 8017 2461
rect 8045 2436 8047 2461
rect 8089 2436 8091 2461
rect 8134 2436 8136 2461
rect 8001 2267 8003 2292
rect 8009 2267 8011 2292
rect 8039 2267 8041 2292
rect 8083 2267 8085 2292
rect 8128 2267 8130 2292
rect 12498 2227 12500 2239
rect 12537 2211 12539 2235
rect 12547 2211 12549 2235
rect 12565 2205 12567 2229
rect 12575 2205 12577 2229
rect 12498 2172 12500 2184
rect 8001 2087 8003 2112
rect 8009 2087 8011 2112
rect 8039 2087 8041 2112
rect 8083 2087 8085 2112
rect 8128 2087 8130 2112
rect 8536 2090 8538 2102
rect 8575 2074 8577 2098
rect 8585 2074 8587 2098
rect 8603 2068 8605 2092
rect 8613 2068 8615 2092
rect 8536 2035 8538 2047
rect 13413 2033 13415 2053
rect 10234 1954 10236 2004
rect 10284 1955 10286 2005
rect 10334 1955 10336 2005
rect 10381 1955 10383 2005
rect 12928 1973 12930 1998
rect 12936 1973 12938 1998
rect 12966 1973 12968 1998
rect 13010 1973 13012 1998
rect 13055 1973 13057 1998
rect 9023 1876 9025 1896
rect 9034 1876 9036 1896
rect 9065 1869 9067 1889
rect 8049 1771 8051 1796
rect 8057 1771 8059 1796
rect 8087 1771 8089 1796
rect 8131 1771 8133 1796
rect 8176 1771 8178 1796
rect 8527 1731 8529 1743
rect 8566 1715 8568 1739
rect 8576 1715 8578 1739
rect 8594 1709 8596 1733
rect 8604 1709 8606 1733
rect 8527 1676 8529 1688
rect 10703 1733 10705 1773
rect 10741 1733 10743 1773
rect 10785 1733 10787 1773
rect 10823 1733 10825 1773
rect 10869 1735 10871 1775
rect 8053 1609 8055 1634
rect 8061 1609 8063 1634
rect 8091 1609 8093 1634
rect 8135 1609 8137 1634
rect 8180 1609 8182 1634
rect 13441 1612 13443 1632
rect 9025 1526 9027 1546
rect 9036 1526 9038 1546
rect 9067 1519 9069 1539
rect 12913 1532 12915 1557
rect 12921 1532 12923 1557
rect 12951 1532 12953 1557
rect 12995 1532 12997 1557
rect 13040 1532 13042 1557
rect 12538 1417 12540 1429
rect 12577 1401 12579 1425
rect 12587 1401 12589 1425
rect 12605 1395 12607 1419
rect 12615 1395 12617 1419
rect 8058 1359 8060 1384
rect 8066 1359 8068 1384
rect 8096 1359 8098 1384
rect 8140 1359 8142 1384
rect 8185 1359 8187 1384
rect 8554 1372 8556 1384
rect 8593 1356 8595 1380
rect 8603 1356 8605 1380
rect 8621 1350 8623 1374
rect 8631 1350 8633 1374
rect 12538 1362 12540 1374
rect 8554 1317 8556 1329
rect 9033 1234 9035 1254
rect 9044 1234 9046 1254
rect 8056 1199 8058 1224
rect 8064 1199 8066 1224
rect 8094 1199 8096 1224
rect 8138 1199 8140 1224
rect 8183 1199 8185 1224
rect 9075 1227 9077 1247
rect 13492 1058 13494 1078
rect 8547 1029 8549 1041
rect 8586 1013 8588 1037
rect 8596 1013 8598 1037
rect 8614 1007 8616 1031
rect 8624 1007 8626 1031
rect 8084 964 8086 989
rect 8092 964 8094 989
rect 8122 964 8124 989
rect 8166 964 8168 989
rect 8211 964 8213 989
rect 8547 974 8549 986
rect 12478 987 12480 999
rect 12517 971 12519 995
rect 12527 971 12529 995
rect 12545 965 12547 989
rect 12555 965 12557 989
rect 12898 979 12900 1004
rect 12906 979 12908 1004
rect 12936 979 12938 1004
rect 12980 979 12982 1004
rect 13025 979 13027 1004
rect 12478 932 12480 944
rect 9021 868 9023 888
rect 9032 868 9034 888
rect 8093 839 8095 864
rect 8101 839 8103 864
rect 8131 839 8133 864
rect 8175 839 8177 864
rect 8220 839 8222 864
rect 9063 861 9065 881
rect 12911 687 12913 712
rect 12919 687 12921 712
rect 12949 687 12951 712
rect 12993 687 12995 712
rect 13038 687 13040 712
rect 13477 709 13479 729
rect 12435 451 12437 463
rect 12474 435 12476 459
rect 12484 435 12486 459
rect 12502 429 12504 453
rect 12512 429 12514 453
rect 12435 396 12437 408
rect 12933 313 12935 338
rect 12941 313 12943 338
rect 12971 313 12973 338
rect 13015 313 13017 338
rect 13060 313 13062 338
rect 13530 324 13532 344
<< ndiffusion >>
rect 8002 2404 8003 2414
rect 8005 2404 8006 2414
rect 8038 2404 8039 2414
rect 8041 2404 8042 2414
rect 8046 2404 8047 2414
rect 8049 2404 8050 2414
rect 8082 2404 8083 2414
rect 8085 2404 8086 2414
rect 8090 2404 8091 2414
rect 8093 2404 8094 2414
rect 8133 2404 8134 2414
rect 8136 2404 8137 2414
rect 7996 2235 7997 2245
rect 7999 2235 8000 2245
rect 8032 2235 8033 2245
rect 8035 2235 8036 2245
rect 8040 2235 8041 2245
rect 8043 2235 8044 2245
rect 8076 2235 8077 2245
rect 8079 2235 8080 2245
rect 8084 2235 8085 2245
rect 8087 2235 8088 2245
rect 8127 2235 8128 2245
rect 8130 2235 8131 2245
rect 12497 2207 12498 2213
rect 12500 2207 12501 2213
rect 12536 2158 12537 2170
rect 12539 2158 12547 2170
rect 12549 2158 12550 2170
rect 12564 2158 12565 2170
rect 12567 2158 12575 2170
rect 12577 2158 12578 2170
rect 12497 2152 12498 2158
rect 12500 2152 12501 2158
rect 8535 2070 8536 2076
rect 8538 2070 8539 2076
rect 7996 2055 7997 2065
rect 7999 2055 8000 2065
rect 8032 2055 8033 2065
rect 8035 2055 8036 2065
rect 8040 2055 8041 2065
rect 8043 2055 8044 2065
rect 8076 2055 8077 2065
rect 8079 2055 8080 2065
rect 8084 2055 8085 2065
rect 8087 2055 8088 2065
rect 8127 2055 8128 2065
rect 8130 2055 8131 2065
rect 8574 2021 8575 2033
rect 8577 2021 8585 2033
rect 8587 2021 8588 2033
rect 8602 2021 8603 2033
rect 8605 2021 8613 2033
rect 8615 2021 8616 2033
rect 8535 2015 8536 2021
rect 8538 2015 8539 2021
rect 13412 2005 13413 2015
rect 13415 2005 13416 2015
rect 12923 1941 12924 1951
rect 12926 1941 12927 1951
rect 12959 1941 12960 1951
rect 12962 1941 12963 1951
rect 12967 1941 12968 1951
rect 12970 1941 12971 1951
rect 13003 1941 13004 1951
rect 13006 1941 13007 1951
rect 13011 1941 13012 1951
rect 13014 1941 13015 1951
rect 13054 1941 13055 1951
rect 13057 1941 13058 1951
rect 9022 1827 9023 1847
rect 9025 1827 9034 1847
rect 9036 1827 9037 1847
rect 9064 1845 9065 1855
rect 9067 1845 9068 1855
rect 8044 1739 8045 1749
rect 8047 1739 8048 1749
rect 8080 1739 8081 1749
rect 8083 1739 8084 1749
rect 8088 1739 8089 1749
rect 8091 1739 8092 1749
rect 8124 1739 8125 1749
rect 8127 1739 8128 1749
rect 8132 1739 8133 1749
rect 8135 1739 8136 1749
rect 8175 1739 8176 1749
rect 8178 1739 8179 1749
rect 8526 1711 8527 1717
rect 8529 1711 8530 1717
rect 8565 1662 8566 1674
rect 8568 1662 8576 1674
rect 8578 1662 8579 1674
rect 8593 1662 8594 1674
rect 8596 1662 8604 1674
rect 8606 1662 8607 1674
rect 10169 1668 10170 1768
rect 10172 1668 10173 1768
rect 10197 1668 10198 1768
rect 10200 1668 10201 1768
rect 10224 1668 10225 1768
rect 10227 1668 10228 1768
rect 10263 1668 10264 1768
rect 10266 1668 10267 1768
rect 10291 1668 10292 1768
rect 10294 1668 10295 1768
rect 10318 1668 10319 1768
rect 10321 1668 10322 1768
rect 10358 1669 10359 1769
rect 10361 1669 10362 1769
rect 10386 1669 10387 1769
rect 10389 1669 10390 1769
rect 10413 1669 10414 1769
rect 10416 1669 10417 1769
rect 10449 1669 10450 1769
rect 10452 1669 10453 1769
rect 10702 1695 10703 1715
rect 10705 1695 10706 1715
rect 10740 1695 10741 1715
rect 10743 1695 10744 1715
rect 10784 1695 10785 1715
rect 10787 1695 10788 1715
rect 10822 1695 10823 1715
rect 10825 1695 10826 1715
rect 10868 1697 10869 1717
rect 10871 1697 10872 1717
rect 8526 1656 8527 1662
rect 8529 1656 8530 1662
rect 8048 1577 8049 1587
rect 8051 1577 8052 1587
rect 8084 1577 8085 1587
rect 8087 1577 8088 1587
rect 8092 1577 8093 1587
rect 8095 1577 8096 1587
rect 8128 1577 8129 1587
rect 8131 1577 8132 1587
rect 8136 1577 8137 1587
rect 8139 1577 8140 1587
rect 8179 1577 8180 1587
rect 8182 1577 8183 1587
rect 13440 1584 13441 1594
rect 13443 1584 13444 1594
rect 9024 1477 9025 1497
rect 9027 1477 9036 1497
rect 9038 1477 9039 1497
rect 9066 1495 9067 1505
rect 9069 1495 9070 1505
rect 12908 1500 12909 1510
rect 12911 1500 12912 1510
rect 12944 1500 12945 1510
rect 12947 1500 12948 1510
rect 12952 1500 12953 1510
rect 12955 1500 12956 1510
rect 12988 1500 12989 1510
rect 12991 1500 12992 1510
rect 12996 1500 12997 1510
rect 12999 1500 13000 1510
rect 13039 1500 13040 1510
rect 13042 1500 13043 1510
rect 12537 1397 12538 1403
rect 12540 1397 12541 1403
rect 8553 1352 8554 1358
rect 8556 1352 8557 1358
rect 8053 1327 8054 1337
rect 8056 1327 8057 1337
rect 8089 1327 8090 1337
rect 8092 1327 8093 1337
rect 8097 1327 8098 1337
rect 8100 1327 8101 1337
rect 8133 1327 8134 1337
rect 8136 1327 8137 1337
rect 8141 1327 8142 1337
rect 8144 1327 8145 1337
rect 8184 1327 8185 1337
rect 8187 1327 8188 1337
rect 12576 1348 12577 1360
rect 12579 1348 12587 1360
rect 12589 1348 12590 1360
rect 12604 1348 12605 1360
rect 12607 1348 12615 1360
rect 12617 1348 12618 1360
rect 12537 1342 12538 1348
rect 12540 1342 12541 1348
rect 8592 1303 8593 1315
rect 8595 1303 8603 1315
rect 8605 1303 8606 1315
rect 8620 1303 8621 1315
rect 8623 1303 8631 1315
rect 8633 1303 8634 1315
rect 8553 1297 8554 1303
rect 8556 1297 8557 1303
rect 9032 1185 9033 1205
rect 9035 1185 9044 1205
rect 9046 1185 9047 1205
rect 9074 1203 9075 1213
rect 9077 1203 9078 1213
rect 8051 1167 8052 1177
rect 8054 1167 8055 1177
rect 8087 1167 8088 1177
rect 8090 1167 8091 1177
rect 8095 1167 8096 1177
rect 8098 1167 8099 1177
rect 8131 1167 8132 1177
rect 8134 1167 8135 1177
rect 8139 1167 8140 1177
rect 8142 1167 8143 1177
rect 8182 1167 8183 1177
rect 8185 1167 8186 1177
rect 8546 1009 8547 1015
rect 8549 1009 8550 1015
rect 13491 1030 13492 1040
rect 13494 1030 13495 1040
rect 8585 960 8586 972
rect 8588 960 8596 972
rect 8598 960 8599 972
rect 8613 960 8614 972
rect 8616 960 8624 972
rect 8626 960 8627 972
rect 12477 967 12478 973
rect 12480 967 12481 973
rect 8546 954 8547 960
rect 8549 954 8550 960
rect 8079 932 8080 942
rect 8082 932 8083 942
rect 8115 932 8116 942
rect 8118 932 8119 942
rect 8123 932 8124 942
rect 8126 932 8127 942
rect 8159 932 8160 942
rect 8162 932 8163 942
rect 8167 932 8168 942
rect 8170 932 8171 942
rect 8210 932 8211 942
rect 8213 932 8214 942
rect 12893 947 12894 957
rect 12896 947 12897 957
rect 12929 947 12930 957
rect 12932 947 12933 957
rect 12937 947 12938 957
rect 12940 947 12941 957
rect 12973 947 12974 957
rect 12976 947 12977 957
rect 12981 947 12982 957
rect 12984 947 12985 957
rect 13024 947 13025 957
rect 13027 947 13028 957
rect 12516 918 12517 930
rect 12519 918 12527 930
rect 12529 918 12530 930
rect 12544 918 12545 930
rect 12547 918 12555 930
rect 12557 918 12558 930
rect 12477 912 12478 918
rect 12480 912 12481 918
rect 9020 819 9021 839
rect 9023 819 9032 839
rect 9034 819 9035 839
rect 9062 837 9063 847
rect 9065 837 9066 847
rect 8088 807 8089 817
rect 8091 807 8092 817
rect 8124 807 8125 817
rect 8127 807 8128 817
rect 8132 807 8133 817
rect 8135 807 8136 817
rect 8168 807 8169 817
rect 8171 807 8172 817
rect 8176 807 8177 817
rect 8179 807 8180 817
rect 8219 807 8220 817
rect 8222 807 8223 817
rect 13476 681 13477 691
rect 13479 681 13480 691
rect 12906 655 12907 665
rect 12909 655 12910 665
rect 12942 655 12943 665
rect 12945 655 12946 665
rect 12950 655 12951 665
rect 12953 655 12954 665
rect 12986 655 12987 665
rect 12989 655 12990 665
rect 12994 655 12995 665
rect 12997 655 12998 665
rect 13037 655 13038 665
rect 13040 655 13041 665
rect 12434 431 12435 437
rect 12437 431 12438 437
rect 12473 382 12474 394
rect 12476 382 12484 394
rect 12486 382 12487 394
rect 12501 382 12502 394
rect 12504 382 12512 394
rect 12514 382 12515 394
rect 12434 376 12435 382
rect 12437 376 12438 382
rect 13529 296 13530 306
rect 13532 296 13533 306
rect 12928 281 12929 291
rect 12931 281 12932 291
rect 12964 281 12965 291
rect 12967 281 12968 291
rect 12972 281 12973 291
rect 12975 281 12976 291
rect 13008 281 13009 291
rect 13011 281 13012 291
rect 13016 281 13017 291
rect 13019 281 13020 291
rect 13059 281 13060 291
rect 13062 281 13063 291
<< pdiffusion >>
rect 8006 2436 8007 2461
rect 8009 2436 8010 2461
rect 8014 2436 8015 2461
rect 8017 2436 8018 2461
rect 8044 2436 8045 2461
rect 8047 2436 8048 2461
rect 8088 2436 8089 2461
rect 8091 2436 8092 2461
rect 8133 2436 8134 2461
rect 8136 2436 8137 2461
rect 8000 2267 8001 2292
rect 8003 2267 8004 2292
rect 8008 2267 8009 2292
rect 8011 2267 8012 2292
rect 8038 2267 8039 2292
rect 8041 2267 8042 2292
rect 8082 2267 8083 2292
rect 8085 2267 8086 2292
rect 8127 2267 8128 2292
rect 8130 2267 8131 2292
rect 12497 2227 12498 2239
rect 12500 2227 12501 2239
rect 12536 2211 12537 2235
rect 12539 2211 12541 2235
rect 12545 2211 12547 2235
rect 12549 2211 12550 2235
rect 12564 2205 12565 2229
rect 12567 2205 12569 2229
rect 12573 2205 12575 2229
rect 12577 2205 12578 2229
rect 12497 2172 12498 2184
rect 12500 2172 12501 2184
rect 8000 2087 8001 2112
rect 8003 2087 8004 2112
rect 8008 2087 8009 2112
rect 8011 2087 8012 2112
rect 8038 2087 8039 2112
rect 8041 2087 8042 2112
rect 8082 2087 8083 2112
rect 8085 2087 8086 2112
rect 8127 2087 8128 2112
rect 8130 2087 8131 2112
rect 8535 2090 8536 2102
rect 8538 2090 8539 2102
rect 8574 2074 8575 2098
rect 8577 2074 8579 2098
rect 8583 2074 8585 2098
rect 8587 2074 8588 2098
rect 8602 2068 8603 2092
rect 8605 2068 8607 2092
rect 8611 2068 8613 2092
rect 8615 2068 8616 2092
rect 8535 2035 8536 2047
rect 8538 2035 8539 2047
rect 13412 2033 13413 2053
rect 13415 2033 13416 2053
rect 10233 1954 10234 2004
rect 10236 1954 10237 2004
rect 10283 1955 10284 2005
rect 10286 1955 10287 2005
rect 10333 1955 10334 2005
rect 10336 1955 10337 2005
rect 10380 1955 10381 2005
rect 10383 1955 10384 2005
rect 12927 1973 12928 1998
rect 12930 1973 12931 1998
rect 12935 1973 12936 1998
rect 12938 1973 12939 1998
rect 12965 1973 12966 1998
rect 12968 1973 12969 1998
rect 13009 1973 13010 1998
rect 13012 1973 13013 1998
rect 13054 1973 13055 1998
rect 13057 1973 13058 1998
rect 9022 1876 9023 1896
rect 9025 1876 9029 1896
rect 9033 1876 9034 1896
rect 9036 1876 9037 1896
rect 9064 1869 9065 1889
rect 9067 1869 9068 1889
rect 8048 1771 8049 1796
rect 8051 1771 8052 1796
rect 8056 1771 8057 1796
rect 8059 1771 8060 1796
rect 8086 1771 8087 1796
rect 8089 1771 8090 1796
rect 8130 1771 8131 1796
rect 8133 1771 8134 1796
rect 8175 1771 8176 1796
rect 8178 1771 8179 1796
rect 8526 1731 8527 1743
rect 8529 1731 8530 1743
rect 8565 1715 8566 1739
rect 8568 1715 8570 1739
rect 8574 1715 8576 1739
rect 8578 1715 8579 1739
rect 8593 1709 8594 1733
rect 8596 1709 8598 1733
rect 8602 1709 8604 1733
rect 8606 1709 8607 1733
rect 8526 1676 8527 1688
rect 8529 1676 8530 1688
rect 10702 1733 10703 1773
rect 10705 1733 10706 1773
rect 10740 1733 10741 1773
rect 10743 1733 10744 1773
rect 10784 1733 10785 1773
rect 10787 1733 10788 1773
rect 10822 1733 10823 1773
rect 10825 1733 10826 1773
rect 10868 1735 10869 1775
rect 10871 1735 10872 1775
rect 8052 1609 8053 1634
rect 8055 1609 8056 1634
rect 8060 1609 8061 1634
rect 8063 1609 8064 1634
rect 8090 1609 8091 1634
rect 8093 1609 8094 1634
rect 8134 1609 8135 1634
rect 8137 1609 8138 1634
rect 8179 1609 8180 1634
rect 8182 1609 8183 1634
rect 13440 1612 13441 1632
rect 13443 1612 13444 1632
rect 9024 1526 9025 1546
rect 9027 1526 9031 1546
rect 9035 1526 9036 1546
rect 9038 1526 9039 1546
rect 9066 1519 9067 1539
rect 9069 1519 9070 1539
rect 12912 1532 12913 1557
rect 12915 1532 12916 1557
rect 12920 1532 12921 1557
rect 12923 1532 12924 1557
rect 12950 1532 12951 1557
rect 12953 1532 12954 1557
rect 12994 1532 12995 1557
rect 12997 1532 12998 1557
rect 13039 1532 13040 1557
rect 13042 1532 13043 1557
rect 12537 1417 12538 1429
rect 12540 1417 12541 1429
rect 12576 1401 12577 1425
rect 12579 1401 12581 1425
rect 12585 1401 12587 1425
rect 12589 1401 12590 1425
rect 12604 1395 12605 1419
rect 12607 1395 12609 1419
rect 12613 1395 12615 1419
rect 12617 1395 12618 1419
rect 8057 1359 8058 1384
rect 8060 1359 8061 1384
rect 8065 1359 8066 1384
rect 8068 1359 8069 1384
rect 8095 1359 8096 1384
rect 8098 1359 8099 1384
rect 8139 1359 8140 1384
rect 8142 1359 8143 1384
rect 8184 1359 8185 1384
rect 8187 1359 8188 1384
rect 8553 1372 8554 1384
rect 8556 1372 8557 1384
rect 8592 1356 8593 1380
rect 8595 1356 8597 1380
rect 8601 1356 8603 1380
rect 8605 1356 8606 1380
rect 8620 1350 8621 1374
rect 8623 1350 8625 1374
rect 8629 1350 8631 1374
rect 8633 1350 8634 1374
rect 12537 1362 12538 1374
rect 12540 1362 12541 1374
rect 8553 1317 8554 1329
rect 8556 1317 8557 1329
rect 9032 1234 9033 1254
rect 9035 1234 9039 1254
rect 9043 1234 9044 1254
rect 9046 1234 9047 1254
rect 8055 1199 8056 1224
rect 8058 1199 8059 1224
rect 8063 1199 8064 1224
rect 8066 1199 8067 1224
rect 8093 1199 8094 1224
rect 8096 1199 8097 1224
rect 8137 1199 8138 1224
rect 8140 1199 8141 1224
rect 8182 1199 8183 1224
rect 8185 1199 8186 1224
rect 9074 1227 9075 1247
rect 9077 1227 9078 1247
rect 13491 1058 13492 1078
rect 13494 1058 13495 1078
rect 8546 1029 8547 1041
rect 8549 1029 8550 1041
rect 8585 1013 8586 1037
rect 8588 1013 8590 1037
rect 8594 1013 8596 1037
rect 8598 1013 8599 1037
rect 8613 1007 8614 1031
rect 8616 1007 8618 1031
rect 8622 1007 8624 1031
rect 8626 1007 8627 1031
rect 8083 964 8084 989
rect 8086 964 8087 989
rect 8091 964 8092 989
rect 8094 964 8095 989
rect 8121 964 8122 989
rect 8124 964 8125 989
rect 8165 964 8166 989
rect 8168 964 8169 989
rect 8210 964 8211 989
rect 8213 964 8214 989
rect 8546 974 8547 986
rect 8549 974 8550 986
rect 12477 987 12478 999
rect 12480 987 12481 999
rect 12516 971 12517 995
rect 12519 971 12521 995
rect 12525 971 12527 995
rect 12529 971 12530 995
rect 12544 965 12545 989
rect 12547 965 12549 989
rect 12553 965 12555 989
rect 12557 965 12558 989
rect 12897 979 12898 1004
rect 12900 979 12901 1004
rect 12905 979 12906 1004
rect 12908 979 12909 1004
rect 12935 979 12936 1004
rect 12938 979 12939 1004
rect 12979 979 12980 1004
rect 12982 979 12983 1004
rect 13024 979 13025 1004
rect 13027 979 13028 1004
rect 12477 932 12478 944
rect 12480 932 12481 944
rect 9020 868 9021 888
rect 9023 868 9027 888
rect 9031 868 9032 888
rect 9034 868 9035 888
rect 8092 839 8093 864
rect 8095 839 8096 864
rect 8100 839 8101 864
rect 8103 839 8104 864
rect 8130 839 8131 864
rect 8133 839 8134 864
rect 8174 839 8175 864
rect 8177 839 8178 864
rect 8219 839 8220 864
rect 8222 839 8223 864
rect 9062 861 9063 881
rect 9065 861 9066 881
rect 12910 687 12911 712
rect 12913 687 12914 712
rect 12918 687 12919 712
rect 12921 687 12922 712
rect 12948 687 12949 712
rect 12951 687 12952 712
rect 12992 687 12993 712
rect 12995 687 12996 712
rect 13037 687 13038 712
rect 13040 687 13041 712
rect 13476 709 13477 729
rect 13479 709 13480 729
rect 12434 451 12435 463
rect 12437 451 12438 463
rect 12473 435 12474 459
rect 12476 435 12478 459
rect 12482 435 12484 459
rect 12486 435 12487 459
rect 12501 429 12502 453
rect 12504 429 12506 453
rect 12510 429 12512 453
rect 12514 429 12515 453
rect 12434 396 12435 408
rect 12437 396 12438 408
rect 12932 313 12933 338
rect 12935 313 12936 338
rect 12940 313 12941 338
rect 12943 313 12944 338
rect 12970 313 12971 338
rect 12973 313 12974 338
rect 13014 313 13015 338
rect 13017 313 13018 338
rect 13059 313 13060 338
rect 13062 313 13063 338
rect 13529 324 13530 344
rect 13532 324 13533 344
<< ndcontact >>
rect 7998 2404 8002 2414
rect 8006 2404 8010 2414
rect 8034 2404 8038 2414
rect 8042 2404 8046 2414
rect 8050 2404 8054 2414
rect 8078 2404 8082 2414
rect 8086 2404 8090 2414
rect 8094 2404 8098 2414
rect 8129 2404 8133 2414
rect 8137 2404 8141 2414
rect 7992 2235 7996 2245
rect 8000 2235 8004 2245
rect 8028 2235 8032 2245
rect 8036 2235 8040 2245
rect 8044 2235 8048 2245
rect 8072 2235 8076 2245
rect 8080 2235 8084 2245
rect 8088 2235 8092 2245
rect 8123 2235 8127 2245
rect 8131 2235 8135 2245
rect 12493 2207 12497 2213
rect 12501 2207 12505 2213
rect 12532 2158 12536 2170
rect 12550 2158 12554 2170
rect 12560 2158 12564 2170
rect 12578 2158 12582 2170
rect 12493 2152 12497 2158
rect 12501 2152 12505 2158
rect 8531 2070 8535 2076
rect 8539 2070 8543 2076
rect 7992 2055 7996 2065
rect 8000 2055 8004 2065
rect 8028 2055 8032 2065
rect 8036 2055 8040 2065
rect 8044 2055 8048 2065
rect 8072 2055 8076 2065
rect 8080 2055 8084 2065
rect 8088 2055 8092 2065
rect 8123 2055 8127 2065
rect 8131 2055 8135 2065
rect 8570 2021 8574 2033
rect 8588 2021 8592 2033
rect 8598 2021 8602 2033
rect 8616 2021 8620 2033
rect 8531 2015 8535 2021
rect 8539 2015 8543 2021
rect 13408 2005 13412 2015
rect 13416 2005 13420 2015
rect 12919 1941 12923 1951
rect 12927 1941 12931 1951
rect 12955 1941 12959 1951
rect 12963 1941 12967 1951
rect 12971 1941 12975 1951
rect 12999 1941 13003 1951
rect 13007 1941 13011 1951
rect 13015 1941 13019 1951
rect 13050 1941 13054 1951
rect 13058 1941 13062 1951
rect 9018 1827 9022 1847
rect 9037 1827 9041 1847
rect 9060 1845 9064 1855
rect 9068 1845 9072 1855
rect 8040 1739 8044 1749
rect 8048 1739 8052 1749
rect 8076 1739 8080 1749
rect 8084 1739 8088 1749
rect 8092 1739 8096 1749
rect 8120 1739 8124 1749
rect 8128 1739 8132 1749
rect 8136 1739 8140 1749
rect 8171 1739 8175 1749
rect 8179 1739 8183 1749
rect 8522 1711 8526 1717
rect 8530 1711 8534 1717
rect 8561 1662 8565 1674
rect 8579 1662 8583 1674
rect 8589 1662 8593 1674
rect 8607 1662 8611 1674
rect 10165 1668 10169 1768
rect 10173 1668 10177 1768
rect 10193 1668 10197 1768
rect 10201 1668 10205 1768
rect 10220 1668 10224 1768
rect 10228 1668 10232 1768
rect 10259 1668 10263 1768
rect 10267 1668 10271 1768
rect 10287 1668 10291 1768
rect 10295 1668 10299 1768
rect 10314 1668 10318 1768
rect 10322 1668 10326 1768
rect 10354 1669 10358 1769
rect 10362 1669 10366 1769
rect 10382 1669 10386 1769
rect 10390 1669 10394 1769
rect 10409 1669 10413 1769
rect 10417 1669 10421 1769
rect 10445 1669 10449 1769
rect 10453 1669 10457 1769
rect 10698 1695 10702 1715
rect 10706 1695 10710 1715
rect 10736 1695 10740 1715
rect 10744 1695 10748 1715
rect 10780 1695 10784 1715
rect 10788 1695 10792 1715
rect 10818 1695 10822 1715
rect 10826 1695 10830 1715
rect 10864 1697 10868 1717
rect 10872 1697 10876 1717
rect 8522 1656 8526 1662
rect 8530 1656 8534 1662
rect 8044 1577 8048 1587
rect 8052 1577 8056 1587
rect 8080 1577 8084 1587
rect 8088 1577 8092 1587
rect 8096 1577 8100 1587
rect 8124 1577 8128 1587
rect 8132 1577 8136 1587
rect 8140 1577 8144 1587
rect 8175 1577 8179 1587
rect 8183 1577 8187 1587
rect 13436 1584 13440 1594
rect 13444 1584 13448 1594
rect 9020 1477 9024 1497
rect 9039 1477 9043 1497
rect 9062 1495 9066 1505
rect 9070 1495 9074 1505
rect 12904 1500 12908 1510
rect 12912 1500 12916 1510
rect 12940 1500 12944 1510
rect 12948 1500 12952 1510
rect 12956 1500 12960 1510
rect 12984 1500 12988 1510
rect 12992 1500 12996 1510
rect 13000 1500 13004 1510
rect 13035 1500 13039 1510
rect 13043 1500 13047 1510
rect 12533 1397 12537 1403
rect 12541 1397 12545 1403
rect 8549 1352 8553 1358
rect 8557 1352 8561 1358
rect 8049 1327 8053 1337
rect 8057 1327 8061 1337
rect 8085 1327 8089 1337
rect 8093 1327 8097 1337
rect 8101 1327 8105 1337
rect 8129 1327 8133 1337
rect 8137 1327 8141 1337
rect 8145 1327 8149 1337
rect 8180 1327 8184 1337
rect 8188 1327 8192 1337
rect 12572 1348 12576 1360
rect 12590 1348 12594 1360
rect 12600 1348 12604 1360
rect 12618 1348 12622 1360
rect 12533 1342 12537 1348
rect 12541 1342 12545 1348
rect 8588 1303 8592 1315
rect 8606 1303 8610 1315
rect 8616 1303 8620 1315
rect 8634 1303 8638 1315
rect 8549 1297 8553 1303
rect 8557 1297 8561 1303
rect 9028 1185 9032 1205
rect 9047 1185 9051 1205
rect 9070 1203 9074 1213
rect 9078 1203 9082 1213
rect 8047 1167 8051 1177
rect 8055 1167 8059 1177
rect 8083 1167 8087 1177
rect 8091 1167 8095 1177
rect 8099 1167 8103 1177
rect 8127 1167 8131 1177
rect 8135 1167 8139 1177
rect 8143 1167 8147 1177
rect 8178 1167 8182 1177
rect 8186 1167 8190 1177
rect 8542 1009 8546 1015
rect 8550 1009 8554 1015
rect 13487 1030 13491 1040
rect 13495 1030 13499 1040
rect 8581 960 8585 972
rect 8599 960 8603 972
rect 8609 960 8613 972
rect 8627 960 8631 972
rect 12473 967 12477 973
rect 12481 967 12485 973
rect 8542 954 8546 960
rect 8550 954 8554 960
rect 8075 932 8079 942
rect 8083 932 8087 942
rect 8111 932 8115 942
rect 8119 932 8123 942
rect 8127 932 8131 942
rect 8155 932 8159 942
rect 8163 932 8167 942
rect 8171 932 8175 942
rect 8206 932 8210 942
rect 8214 932 8218 942
rect 12889 947 12893 957
rect 12897 947 12901 957
rect 12925 947 12929 957
rect 12933 947 12937 957
rect 12941 947 12945 957
rect 12969 947 12973 957
rect 12977 947 12981 957
rect 12985 947 12989 957
rect 13020 947 13024 957
rect 13028 947 13032 957
rect 12512 918 12516 930
rect 12530 918 12534 930
rect 12540 918 12544 930
rect 12558 918 12562 930
rect 12473 912 12477 918
rect 12481 912 12485 918
rect 9016 819 9020 839
rect 9035 819 9039 839
rect 9058 837 9062 847
rect 9066 837 9070 847
rect 8084 807 8088 817
rect 8092 807 8096 817
rect 8120 807 8124 817
rect 8128 807 8132 817
rect 8136 807 8140 817
rect 8164 807 8168 817
rect 8172 807 8176 817
rect 8180 807 8184 817
rect 8215 807 8219 817
rect 8223 807 8227 817
rect 13472 681 13476 691
rect 13480 681 13484 691
rect 12902 655 12906 665
rect 12910 655 12914 665
rect 12938 655 12942 665
rect 12946 655 12950 665
rect 12954 655 12958 665
rect 12982 655 12986 665
rect 12990 655 12994 665
rect 12998 655 13002 665
rect 13033 655 13037 665
rect 13041 655 13045 665
rect 12430 431 12434 437
rect 12438 431 12442 437
rect 12469 382 12473 394
rect 12487 382 12491 394
rect 12497 382 12501 394
rect 12515 382 12519 394
rect 12430 376 12434 382
rect 12438 376 12442 382
rect 13525 296 13529 306
rect 13533 296 13537 306
rect 12924 281 12928 291
rect 12932 281 12936 291
rect 12960 281 12964 291
rect 12968 281 12972 291
rect 12976 281 12980 291
rect 13004 281 13008 291
rect 13012 281 13016 291
rect 13020 281 13024 291
rect 13055 281 13059 291
rect 13063 281 13067 291
<< pdcontact >>
rect 8002 2436 8006 2461
rect 8010 2436 8014 2461
rect 8018 2436 8022 2461
rect 8040 2436 8044 2461
rect 8048 2436 8052 2461
rect 8084 2436 8088 2461
rect 8092 2436 8096 2461
rect 8129 2436 8133 2461
rect 8137 2436 8141 2461
rect 7996 2267 8000 2292
rect 8004 2267 8008 2292
rect 8012 2267 8016 2292
rect 8034 2267 8038 2292
rect 8042 2267 8046 2292
rect 8078 2267 8082 2292
rect 8086 2267 8090 2292
rect 8123 2267 8127 2292
rect 8131 2267 8135 2292
rect 12493 2227 12497 2239
rect 12501 2227 12505 2239
rect 12532 2211 12536 2235
rect 12541 2211 12545 2235
rect 12550 2211 12554 2235
rect 12560 2205 12564 2229
rect 12569 2205 12573 2229
rect 12578 2205 12582 2229
rect 12493 2172 12497 2184
rect 12501 2172 12505 2184
rect 7996 2087 8000 2112
rect 8004 2087 8008 2112
rect 8012 2087 8016 2112
rect 8034 2087 8038 2112
rect 8042 2087 8046 2112
rect 8078 2087 8082 2112
rect 8086 2087 8090 2112
rect 8123 2087 8127 2112
rect 8131 2087 8135 2112
rect 8531 2090 8535 2102
rect 8539 2090 8543 2102
rect 8570 2074 8574 2098
rect 8579 2074 8583 2098
rect 8588 2074 8592 2098
rect 8598 2068 8602 2092
rect 8607 2068 8611 2092
rect 8616 2068 8620 2092
rect 8531 2035 8535 2047
rect 8539 2035 8543 2047
rect 13408 2033 13412 2053
rect 13416 2033 13420 2053
rect 10229 1954 10233 2004
rect 10237 1954 10241 2004
rect 10279 1955 10283 2005
rect 10287 1955 10291 2005
rect 10329 1955 10333 2005
rect 10337 1955 10341 2005
rect 10376 1955 10380 2005
rect 10384 1955 10388 2005
rect 12923 1973 12927 1998
rect 12931 1973 12935 1998
rect 12939 1973 12943 1998
rect 12961 1973 12965 1998
rect 12969 1973 12973 1998
rect 13005 1973 13009 1998
rect 13013 1973 13017 1998
rect 13050 1973 13054 1998
rect 13058 1973 13062 1998
rect 9018 1876 9022 1896
rect 9029 1876 9033 1896
rect 9037 1876 9041 1896
rect 9060 1869 9064 1889
rect 9068 1869 9072 1889
rect 8044 1771 8048 1796
rect 8052 1771 8056 1796
rect 8060 1771 8064 1796
rect 8082 1771 8086 1796
rect 8090 1771 8094 1796
rect 8126 1771 8130 1796
rect 8134 1771 8138 1796
rect 8171 1771 8175 1796
rect 8179 1771 8183 1796
rect 8522 1731 8526 1743
rect 8530 1731 8534 1743
rect 8561 1715 8565 1739
rect 8570 1715 8574 1739
rect 8579 1715 8583 1739
rect 8589 1709 8593 1733
rect 8598 1709 8602 1733
rect 8607 1709 8611 1733
rect 8522 1676 8526 1688
rect 8530 1676 8534 1688
rect 10698 1733 10702 1773
rect 10706 1733 10710 1773
rect 10736 1733 10740 1773
rect 10744 1733 10748 1773
rect 10780 1733 10784 1773
rect 10788 1733 10792 1773
rect 10818 1733 10822 1773
rect 10826 1733 10830 1773
rect 10864 1735 10868 1775
rect 10872 1735 10876 1775
rect 8048 1609 8052 1634
rect 8056 1609 8060 1634
rect 8064 1609 8068 1634
rect 8086 1609 8090 1634
rect 8094 1609 8098 1634
rect 8130 1609 8134 1634
rect 8138 1609 8142 1634
rect 8175 1609 8179 1634
rect 8183 1609 8187 1634
rect 13436 1612 13440 1632
rect 13444 1612 13448 1632
rect 9020 1526 9024 1546
rect 9031 1526 9035 1546
rect 9039 1526 9043 1546
rect 9062 1519 9066 1539
rect 9070 1519 9074 1539
rect 12908 1532 12912 1557
rect 12916 1532 12920 1557
rect 12924 1532 12928 1557
rect 12946 1532 12950 1557
rect 12954 1532 12958 1557
rect 12990 1532 12994 1557
rect 12998 1532 13002 1557
rect 13035 1532 13039 1557
rect 13043 1532 13047 1557
rect 12533 1417 12537 1429
rect 12541 1417 12545 1429
rect 12572 1401 12576 1425
rect 12581 1401 12585 1425
rect 12590 1401 12594 1425
rect 12600 1395 12604 1419
rect 12609 1395 12613 1419
rect 12618 1395 12622 1419
rect 8053 1359 8057 1384
rect 8061 1359 8065 1384
rect 8069 1359 8073 1384
rect 8091 1359 8095 1384
rect 8099 1359 8103 1384
rect 8135 1359 8139 1384
rect 8143 1359 8147 1384
rect 8180 1359 8184 1384
rect 8188 1359 8192 1384
rect 8549 1372 8553 1384
rect 8557 1372 8561 1384
rect 8588 1356 8592 1380
rect 8597 1356 8601 1380
rect 8606 1356 8610 1380
rect 8616 1350 8620 1374
rect 8625 1350 8629 1374
rect 8634 1350 8638 1374
rect 12533 1362 12537 1374
rect 12541 1362 12545 1374
rect 8549 1317 8553 1329
rect 8557 1317 8561 1329
rect 9028 1234 9032 1254
rect 9039 1234 9043 1254
rect 9047 1234 9051 1254
rect 8051 1199 8055 1224
rect 8059 1199 8063 1224
rect 8067 1199 8071 1224
rect 8089 1199 8093 1224
rect 8097 1199 8101 1224
rect 8133 1199 8137 1224
rect 8141 1199 8145 1224
rect 8178 1199 8182 1224
rect 8186 1199 8190 1224
rect 9070 1227 9074 1247
rect 9078 1227 9082 1247
rect 13487 1058 13491 1078
rect 13495 1058 13499 1078
rect 8542 1029 8546 1041
rect 8550 1029 8554 1041
rect 8581 1013 8585 1037
rect 8590 1013 8594 1037
rect 8599 1013 8603 1037
rect 8609 1007 8613 1031
rect 8618 1007 8622 1031
rect 8627 1007 8631 1031
rect 8079 964 8083 989
rect 8087 964 8091 989
rect 8095 964 8099 989
rect 8117 964 8121 989
rect 8125 964 8129 989
rect 8161 964 8165 989
rect 8169 964 8173 989
rect 8206 964 8210 989
rect 8214 964 8218 989
rect 8542 974 8546 986
rect 8550 974 8554 986
rect 12473 987 12477 999
rect 12481 987 12485 999
rect 12512 971 12516 995
rect 12521 971 12525 995
rect 12530 971 12534 995
rect 12540 965 12544 989
rect 12549 965 12553 989
rect 12558 965 12562 989
rect 12893 979 12897 1004
rect 12901 979 12905 1004
rect 12909 979 12913 1004
rect 12931 979 12935 1004
rect 12939 979 12943 1004
rect 12975 979 12979 1004
rect 12983 979 12987 1004
rect 13020 979 13024 1004
rect 13028 979 13032 1004
rect 12473 932 12477 944
rect 12481 932 12485 944
rect 9016 868 9020 888
rect 9027 868 9031 888
rect 9035 868 9039 888
rect 8088 839 8092 864
rect 8096 839 8100 864
rect 8104 839 8108 864
rect 8126 839 8130 864
rect 8134 839 8138 864
rect 8170 839 8174 864
rect 8178 839 8182 864
rect 8215 839 8219 864
rect 8223 839 8227 864
rect 9058 861 9062 881
rect 9066 861 9070 881
rect 12906 687 12910 712
rect 12914 687 12918 712
rect 12922 687 12926 712
rect 12944 687 12948 712
rect 12952 687 12956 712
rect 12988 687 12992 712
rect 12996 687 13000 712
rect 13033 687 13037 712
rect 13041 687 13045 712
rect 13472 709 13476 729
rect 13480 709 13484 729
rect 12430 451 12434 463
rect 12438 451 12442 463
rect 12469 435 12473 459
rect 12478 435 12482 459
rect 12487 435 12491 459
rect 12497 429 12501 453
rect 12506 429 12510 453
rect 12515 429 12519 453
rect 12430 396 12434 408
rect 12438 396 12442 408
rect 12928 313 12932 338
rect 12936 313 12940 338
rect 12944 313 12948 338
rect 12966 313 12970 338
rect 12974 313 12978 338
rect 13010 313 13014 338
rect 13018 313 13022 338
rect 13055 313 13059 338
rect 13063 313 13067 338
rect 13525 324 13529 344
rect 13533 324 13537 344
<< psubstratepcontact >>
rect 9074 1836 9079 1840
rect 9076 1486 9081 1490
rect 9084 1194 9089 1198
rect 9072 828 9077 832
<< nsubstratencontact >>
rect 13403 2059 13407 2063
rect 10224 2010 10228 2015
rect 10274 2011 10278 2016
rect 10324 2011 10328 2016
rect 10371 2011 10375 2016
rect 9018 1901 9022 1907
rect 9070 1896 9074 1900
rect 10693 1779 10697 1783
rect 10731 1779 10735 1783
rect 10775 1779 10779 1783
rect 10813 1779 10817 1783
rect 10859 1781 10863 1785
rect 13431 1638 13435 1642
rect 9020 1551 9024 1557
rect 9072 1546 9076 1550
rect 9028 1259 9032 1265
rect 9080 1254 9084 1258
rect 13482 1084 13486 1088
rect 9016 893 9020 899
rect 9068 888 9072 892
rect 13467 735 13471 739
rect 13520 350 13524 354
<< polysilicon >>
rect 8007 2461 8009 2464
rect 8015 2461 8017 2464
rect 8045 2461 8047 2464
rect 8089 2461 8091 2464
rect 8134 2461 8136 2464
rect 8007 2429 8009 2436
rect 8002 2425 8009 2429
rect 8003 2414 8005 2425
rect 8015 2417 8017 2436
rect 8045 2428 8047 2436
rect 8089 2428 8091 2436
rect 8039 2426 8047 2428
rect 8083 2426 8091 2428
rect 8039 2414 8041 2426
rect 8047 2414 8049 2423
rect 8083 2414 8085 2426
rect 8091 2414 8093 2423
rect 8134 2414 8136 2436
rect 8003 2401 8005 2404
rect 8039 2401 8041 2404
rect 8047 2401 8049 2404
rect 8083 2401 8085 2404
rect 8091 2401 8093 2404
rect 8134 2401 8136 2404
rect 8001 2292 8003 2295
rect 8009 2292 8011 2295
rect 8039 2292 8041 2295
rect 8083 2292 8085 2295
rect 8128 2292 8130 2295
rect 8001 2260 8003 2267
rect 7996 2256 8003 2260
rect 7997 2245 7999 2256
rect 8009 2248 8011 2267
rect 8039 2259 8041 2267
rect 8083 2259 8085 2267
rect 8033 2257 8041 2259
rect 8077 2257 8085 2259
rect 8033 2245 8035 2257
rect 8041 2245 8043 2254
rect 8077 2245 8079 2257
rect 8085 2245 8087 2254
rect 8128 2245 8130 2267
rect 12498 2239 12500 2242
rect 7997 2232 7999 2235
rect 8033 2232 8035 2235
rect 8041 2232 8043 2235
rect 8077 2232 8079 2235
rect 8085 2232 8087 2235
rect 8128 2232 8130 2235
rect 12537 2235 12539 2238
rect 12547 2235 12549 2238
rect 12498 2213 12500 2227
rect 12565 2229 12567 2232
rect 12575 2229 12577 2232
rect 12498 2204 12500 2207
rect 12537 2202 12539 2211
rect 12547 2201 12549 2211
rect 12498 2184 12500 2187
rect 12498 2158 12500 2172
rect 12537 2170 12539 2197
rect 12547 2170 12549 2196
rect 12565 2194 12567 2205
rect 12565 2170 12567 2190
rect 12575 2183 12577 2205
rect 12575 2170 12577 2179
rect 12537 2155 12539 2158
rect 12547 2155 12549 2158
rect 12565 2155 12567 2158
rect 12575 2155 12577 2158
rect 12498 2149 12500 2152
rect 8001 2112 8003 2115
rect 8009 2112 8011 2115
rect 8039 2112 8041 2115
rect 8083 2112 8085 2115
rect 8128 2112 8130 2115
rect 8536 2102 8538 2105
rect 8575 2098 8577 2101
rect 8585 2098 8587 2101
rect 8001 2080 8003 2087
rect 7996 2076 8003 2080
rect 7997 2065 7999 2076
rect 8009 2068 8011 2087
rect 8039 2079 8041 2087
rect 8083 2079 8085 2087
rect 8033 2077 8041 2079
rect 8077 2077 8085 2079
rect 8033 2065 8035 2077
rect 8041 2065 8043 2074
rect 8077 2065 8079 2077
rect 8085 2065 8087 2074
rect 8128 2065 8130 2087
rect 8536 2076 8538 2090
rect 8603 2092 8605 2095
rect 8613 2092 8615 2095
rect 8536 2067 8538 2070
rect 8575 2065 8577 2074
rect 8585 2064 8587 2074
rect 7997 2052 7999 2055
rect 8033 2052 8035 2055
rect 8041 2052 8043 2055
rect 8077 2052 8079 2055
rect 8085 2052 8087 2055
rect 8128 2052 8130 2055
rect 8536 2047 8538 2050
rect 8536 2021 8538 2035
rect 8575 2033 8577 2060
rect 8585 2033 8587 2059
rect 8603 2057 8605 2068
rect 8603 2033 8605 2053
rect 8613 2046 8615 2068
rect 13413 2053 13415 2056
rect 8613 2033 8615 2042
rect 8575 2018 8577 2021
rect 8585 2018 8587 2021
rect 8603 2018 8605 2021
rect 8613 2018 8615 2021
rect 8536 2012 8538 2015
rect 13413 2015 13415 2033
rect 10234 2004 10236 2007
rect 10284 2005 10286 2008
rect 10334 2005 10336 2008
rect 10381 2005 10383 2008
rect 13413 2001 13415 2005
rect 12928 1998 12930 2001
rect 12936 1998 12938 2001
rect 12966 1998 12968 2001
rect 13010 1998 13012 2001
rect 13055 1998 13057 2001
rect 12928 1966 12930 1973
rect 12923 1962 12930 1966
rect 10234 1931 10236 1954
rect 10284 1932 10286 1955
rect 10334 1932 10336 1955
rect 10381 1932 10383 1955
rect 12924 1951 12926 1962
rect 12936 1954 12938 1973
rect 12966 1965 12968 1973
rect 13010 1965 13012 1973
rect 12960 1963 12968 1965
rect 13004 1963 13012 1965
rect 12960 1951 12962 1963
rect 12968 1951 12970 1960
rect 13004 1951 13006 1963
rect 13012 1951 13014 1960
rect 13055 1951 13057 1973
rect 12924 1938 12926 1941
rect 12960 1938 12962 1941
rect 12968 1938 12970 1941
rect 13004 1938 13006 1941
rect 13012 1938 13014 1941
rect 13055 1938 13057 1941
rect 9023 1896 9025 1899
rect 9034 1896 9036 1899
rect 9065 1889 9067 1893
rect 9023 1847 9025 1876
rect 9034 1847 9036 1876
rect 9065 1855 9067 1869
rect 9065 1842 9067 1845
rect 9023 1824 9025 1827
rect 9034 1824 9036 1827
rect 8049 1796 8051 1799
rect 8057 1796 8059 1799
rect 8087 1796 8089 1799
rect 8131 1796 8133 1799
rect 8176 1796 8178 1799
rect 10703 1773 10705 1776
rect 10741 1773 10743 1776
rect 10785 1773 10787 1776
rect 10823 1773 10825 1776
rect 10869 1775 10871 1778
rect 8049 1764 8051 1771
rect 8044 1760 8051 1764
rect 8045 1749 8047 1760
rect 8057 1752 8059 1771
rect 8087 1763 8089 1771
rect 8131 1763 8133 1771
rect 8081 1761 8089 1763
rect 8125 1761 8133 1763
rect 8081 1749 8083 1761
rect 8089 1749 8091 1758
rect 8125 1749 8127 1761
rect 8133 1749 8135 1758
rect 8176 1749 8178 1771
rect 10170 1768 10172 1771
rect 10198 1768 10200 1771
rect 10225 1768 10227 1771
rect 10264 1768 10266 1771
rect 10292 1768 10294 1771
rect 10319 1768 10321 1771
rect 10359 1769 10361 1772
rect 10387 1769 10389 1772
rect 10414 1769 10416 1772
rect 10450 1769 10452 1772
rect 8527 1743 8529 1746
rect 8045 1736 8047 1739
rect 8081 1736 8083 1739
rect 8089 1736 8091 1739
rect 8125 1736 8127 1739
rect 8133 1736 8135 1739
rect 8176 1736 8178 1739
rect 8566 1739 8568 1742
rect 8576 1739 8578 1742
rect 8527 1717 8529 1731
rect 8594 1733 8596 1736
rect 8604 1733 8606 1736
rect 8527 1708 8529 1711
rect 8566 1706 8568 1715
rect 8576 1705 8578 1715
rect 8527 1688 8529 1691
rect 8527 1662 8529 1676
rect 8566 1674 8568 1701
rect 8576 1674 8578 1700
rect 8594 1698 8596 1709
rect 8594 1674 8596 1694
rect 8604 1687 8606 1709
rect 8604 1674 8606 1683
rect 10703 1715 10705 1733
rect 10741 1715 10743 1733
rect 10785 1715 10787 1733
rect 10823 1715 10825 1733
rect 10869 1717 10871 1735
rect 10703 1691 10705 1695
rect 10741 1691 10743 1695
rect 10785 1691 10787 1695
rect 10823 1691 10825 1695
rect 10869 1693 10871 1697
rect 8566 1659 8568 1662
rect 8576 1659 8578 1662
rect 8594 1659 8596 1662
rect 8604 1659 8606 1662
rect 10170 1656 10172 1668
rect 10198 1656 10200 1668
rect 10225 1656 10227 1668
rect 10264 1656 10266 1668
rect 10292 1656 10294 1668
rect 10319 1656 10321 1668
rect 10359 1657 10361 1669
rect 10387 1657 10389 1669
rect 10414 1657 10416 1669
rect 10450 1657 10452 1669
rect 8527 1653 8529 1656
rect 8053 1634 8055 1637
rect 8061 1634 8063 1637
rect 8091 1634 8093 1637
rect 8135 1634 8137 1637
rect 8180 1634 8182 1637
rect 13441 1632 13443 1635
rect 8053 1602 8055 1609
rect 8048 1598 8055 1602
rect 8049 1587 8051 1598
rect 8061 1590 8063 1609
rect 8091 1601 8093 1609
rect 8135 1601 8137 1609
rect 8085 1599 8093 1601
rect 8129 1599 8137 1601
rect 8085 1587 8087 1599
rect 8093 1587 8095 1596
rect 8129 1587 8131 1599
rect 8137 1587 8139 1596
rect 8180 1587 8182 1609
rect 13441 1594 13443 1612
rect 13441 1580 13443 1584
rect 8049 1574 8051 1577
rect 8085 1574 8087 1577
rect 8093 1574 8095 1577
rect 8129 1574 8131 1577
rect 8137 1574 8139 1577
rect 8180 1574 8182 1577
rect 12913 1557 12915 1560
rect 12921 1557 12923 1560
rect 12951 1557 12953 1560
rect 12995 1557 12997 1560
rect 13040 1557 13042 1560
rect 9025 1546 9027 1549
rect 9036 1546 9038 1549
rect 9067 1539 9069 1543
rect 9025 1497 9027 1526
rect 9036 1497 9038 1526
rect 12913 1525 12915 1532
rect 12908 1521 12915 1525
rect 9067 1505 9069 1519
rect 12909 1510 12911 1521
rect 12921 1513 12923 1532
rect 12951 1524 12953 1532
rect 12995 1524 12997 1532
rect 12945 1522 12953 1524
rect 12989 1522 12997 1524
rect 12945 1510 12947 1522
rect 12953 1510 12955 1519
rect 12989 1510 12991 1522
rect 12997 1510 12999 1519
rect 13040 1510 13042 1532
rect 12909 1497 12911 1500
rect 12945 1497 12947 1500
rect 12953 1497 12955 1500
rect 12989 1497 12991 1500
rect 12997 1497 12999 1500
rect 13040 1497 13042 1500
rect 9067 1492 9069 1495
rect 9025 1474 9027 1477
rect 9036 1474 9038 1477
rect 12538 1429 12540 1432
rect 12577 1425 12579 1428
rect 12587 1425 12589 1428
rect 12538 1403 12540 1417
rect 12605 1419 12607 1422
rect 12615 1419 12617 1422
rect 12538 1394 12540 1397
rect 12577 1392 12579 1401
rect 12587 1391 12589 1401
rect 8058 1384 8060 1387
rect 8066 1384 8068 1387
rect 8096 1384 8098 1387
rect 8140 1384 8142 1387
rect 8185 1384 8187 1387
rect 8554 1384 8556 1387
rect 8593 1380 8595 1383
rect 8603 1380 8605 1383
rect 8058 1352 8060 1359
rect 8053 1348 8060 1352
rect 8054 1337 8056 1348
rect 8066 1340 8068 1359
rect 8096 1351 8098 1359
rect 8140 1351 8142 1359
rect 8090 1349 8098 1351
rect 8134 1349 8142 1351
rect 8090 1337 8092 1349
rect 8098 1337 8100 1346
rect 8134 1337 8136 1349
rect 8142 1337 8144 1346
rect 8185 1337 8187 1359
rect 8554 1358 8556 1372
rect 8621 1374 8623 1377
rect 8631 1374 8633 1377
rect 12538 1374 12540 1377
rect 8554 1349 8556 1352
rect 8593 1347 8595 1356
rect 8603 1346 8605 1356
rect 8554 1329 8556 1332
rect 8054 1324 8056 1327
rect 8090 1324 8092 1327
rect 8098 1324 8100 1327
rect 8134 1324 8136 1327
rect 8142 1324 8144 1327
rect 8185 1324 8187 1327
rect 8554 1303 8556 1317
rect 8593 1315 8595 1342
rect 8603 1315 8605 1341
rect 8621 1339 8623 1350
rect 8621 1315 8623 1335
rect 8631 1328 8633 1350
rect 12538 1348 12540 1362
rect 12577 1360 12579 1387
rect 12587 1360 12589 1386
rect 12605 1384 12607 1395
rect 12605 1360 12607 1380
rect 12615 1373 12617 1395
rect 12615 1360 12617 1369
rect 12577 1345 12579 1348
rect 12587 1345 12589 1348
rect 12605 1345 12607 1348
rect 12615 1345 12617 1348
rect 12538 1339 12540 1342
rect 8631 1315 8633 1324
rect 8593 1300 8595 1303
rect 8603 1300 8605 1303
rect 8621 1300 8623 1303
rect 8631 1300 8633 1303
rect 8554 1294 8556 1297
rect 9033 1254 9035 1257
rect 9044 1254 9046 1257
rect 9075 1247 9077 1251
rect 8056 1224 8058 1227
rect 8064 1224 8066 1227
rect 8094 1224 8096 1227
rect 8138 1224 8140 1227
rect 8183 1224 8185 1227
rect 9033 1205 9035 1234
rect 9044 1205 9046 1234
rect 9075 1213 9077 1227
rect 8056 1192 8058 1199
rect 8051 1188 8058 1192
rect 8052 1177 8054 1188
rect 8064 1180 8066 1199
rect 8094 1191 8096 1199
rect 8138 1191 8140 1199
rect 8088 1189 8096 1191
rect 8132 1189 8140 1191
rect 8088 1177 8090 1189
rect 8096 1177 8098 1186
rect 8132 1177 8134 1189
rect 8140 1177 8142 1186
rect 8183 1177 8185 1199
rect 9075 1200 9077 1203
rect 9033 1182 9035 1185
rect 9044 1182 9046 1185
rect 8052 1164 8054 1167
rect 8088 1164 8090 1167
rect 8096 1164 8098 1167
rect 8132 1164 8134 1167
rect 8140 1164 8142 1167
rect 8183 1164 8185 1167
rect 13492 1078 13494 1081
rect 8547 1041 8549 1044
rect 13492 1040 13494 1058
rect 8586 1037 8588 1040
rect 8596 1037 8598 1040
rect 8547 1015 8549 1029
rect 8614 1031 8616 1034
rect 8624 1031 8626 1034
rect 8547 1006 8549 1009
rect 8586 1004 8588 1013
rect 8596 1003 8598 1013
rect 13492 1026 13494 1030
rect 8084 989 8086 992
rect 8092 989 8094 992
rect 8122 989 8124 992
rect 8166 989 8168 992
rect 8211 989 8213 992
rect 8547 986 8549 989
rect 8084 957 8086 964
rect 8079 953 8086 957
rect 8080 942 8082 953
rect 8092 945 8094 964
rect 8122 956 8124 964
rect 8166 956 8168 964
rect 8116 954 8124 956
rect 8160 954 8168 956
rect 8116 942 8118 954
rect 8124 942 8126 951
rect 8160 942 8162 954
rect 8168 942 8170 951
rect 8211 942 8213 964
rect 8547 960 8549 974
rect 8586 972 8588 999
rect 8596 972 8598 998
rect 8614 996 8616 1007
rect 8614 972 8616 992
rect 8624 985 8626 1007
rect 12898 1004 12900 1007
rect 12906 1004 12908 1007
rect 12936 1004 12938 1007
rect 12980 1004 12982 1007
rect 13025 1004 13027 1007
rect 12478 999 12480 1002
rect 12517 995 12519 998
rect 12527 995 12529 998
rect 8624 972 8626 981
rect 12478 973 12480 987
rect 12545 989 12547 992
rect 12555 989 12557 992
rect 12478 964 12480 967
rect 12517 962 12519 971
rect 8586 957 8588 960
rect 8596 957 8598 960
rect 8614 957 8616 960
rect 8624 957 8626 960
rect 12527 961 12529 971
rect 12898 972 12900 979
rect 12893 968 12900 972
rect 8547 951 8549 954
rect 12478 944 12480 947
rect 8080 929 8082 932
rect 8116 929 8118 932
rect 8124 929 8126 932
rect 8160 929 8162 932
rect 8168 929 8170 932
rect 8211 929 8213 932
rect 12478 918 12480 932
rect 12517 930 12519 957
rect 12527 930 12529 956
rect 12545 954 12547 965
rect 12545 930 12547 950
rect 12555 943 12557 965
rect 12894 957 12896 968
rect 12906 960 12908 979
rect 12936 971 12938 979
rect 12980 971 12982 979
rect 12930 969 12938 971
rect 12974 969 12982 971
rect 12930 957 12932 969
rect 12938 957 12940 966
rect 12974 957 12976 969
rect 12982 957 12984 966
rect 13025 957 13027 979
rect 12894 944 12896 947
rect 12930 944 12932 947
rect 12938 944 12940 947
rect 12974 944 12976 947
rect 12982 944 12984 947
rect 13025 944 13027 947
rect 12555 930 12557 939
rect 12517 915 12519 918
rect 12527 915 12529 918
rect 12545 915 12547 918
rect 12555 915 12557 918
rect 12478 909 12480 912
rect 9021 888 9023 891
rect 9032 888 9034 891
rect 9063 881 9065 885
rect 8093 864 8095 867
rect 8101 864 8103 867
rect 8131 864 8133 867
rect 8175 864 8177 867
rect 8220 864 8222 867
rect 9021 839 9023 868
rect 9032 839 9034 868
rect 9063 847 9065 861
rect 8093 832 8095 839
rect 8088 828 8095 832
rect 8089 817 8091 828
rect 8101 820 8103 839
rect 8131 831 8133 839
rect 8175 831 8177 839
rect 8125 829 8133 831
rect 8169 829 8177 831
rect 8125 817 8127 829
rect 8133 817 8135 826
rect 8169 817 8171 829
rect 8177 817 8179 826
rect 8220 817 8222 839
rect 9063 834 9065 837
rect 9021 816 9023 819
rect 9032 816 9034 819
rect 8089 804 8091 807
rect 8125 804 8127 807
rect 8133 804 8135 807
rect 8169 804 8171 807
rect 8177 804 8179 807
rect 8220 804 8222 807
rect 13477 729 13479 732
rect 12911 712 12913 715
rect 12919 712 12921 715
rect 12949 712 12951 715
rect 12993 712 12995 715
rect 13038 712 13040 715
rect 13477 691 13479 709
rect 12911 680 12913 687
rect 12906 676 12913 680
rect 12907 665 12909 676
rect 12919 668 12921 687
rect 12949 679 12951 687
rect 12993 679 12995 687
rect 12943 677 12951 679
rect 12987 677 12995 679
rect 12943 665 12945 677
rect 12951 665 12953 674
rect 12987 665 12989 677
rect 12995 665 12997 674
rect 13038 665 13040 687
rect 13477 677 13479 681
rect 12907 652 12909 655
rect 12943 652 12945 655
rect 12951 652 12953 655
rect 12987 652 12989 655
rect 12995 652 12997 655
rect 13038 652 13040 655
rect 12435 463 12437 466
rect 12474 459 12476 462
rect 12484 459 12486 462
rect 12435 437 12437 451
rect 12502 453 12504 456
rect 12512 453 12514 456
rect 12435 428 12437 431
rect 12474 426 12476 435
rect 12484 425 12486 435
rect 12435 408 12437 411
rect 12435 382 12437 396
rect 12474 394 12476 421
rect 12484 394 12486 420
rect 12502 418 12504 429
rect 12502 394 12504 414
rect 12512 407 12514 429
rect 12512 394 12514 403
rect 12474 379 12476 382
rect 12484 379 12486 382
rect 12502 379 12504 382
rect 12512 379 12514 382
rect 12435 373 12437 376
rect 13530 344 13532 347
rect 12933 338 12935 341
rect 12941 338 12943 341
rect 12971 338 12973 341
rect 13015 338 13017 341
rect 13060 338 13062 341
rect 12933 306 12935 313
rect 12928 302 12935 306
rect 12929 291 12931 302
rect 12941 294 12943 313
rect 12971 305 12973 313
rect 13015 305 13017 313
rect 12965 303 12973 305
rect 13009 303 13017 305
rect 12965 291 12967 303
rect 12973 291 12975 300
rect 13009 291 13011 303
rect 13017 291 13019 300
rect 13060 291 13062 313
rect 13530 306 13532 324
rect 13530 292 13532 296
rect 12929 278 12931 281
rect 12965 278 12967 281
rect 12973 278 12975 281
rect 13009 278 13011 281
rect 13017 278 13019 281
rect 13060 278 13062 281
<< polycontact >>
rect 7998 2425 8002 2429
rect 8011 2417 8015 2421
rect 8022 2425 8026 2429
rect 8034 2417 8039 2422
rect 8049 2417 8053 2421
rect 8078 2417 8083 2422
rect 8130 2422 8134 2427
rect 8093 2417 8097 2421
rect 7992 2256 7996 2260
rect 8005 2248 8009 2252
rect 8016 2256 8020 2260
rect 8028 2248 8033 2253
rect 8043 2248 8047 2252
rect 8072 2248 8077 2253
rect 8124 2253 8128 2258
rect 8087 2248 8091 2252
rect 12494 2216 12498 2220
rect 12494 2161 12498 2165
rect 12563 2190 12567 2194
rect 12574 2179 12578 2183
rect 7992 2076 7996 2080
rect 8005 2068 8009 2072
rect 8016 2076 8020 2080
rect 8028 2068 8033 2073
rect 8043 2068 8047 2072
rect 8072 2068 8077 2073
rect 8124 2073 8128 2078
rect 8087 2068 8091 2072
rect 8532 2079 8536 2083
rect 8532 2024 8536 2028
rect 8601 2053 8605 2057
rect 8612 2042 8616 2046
rect 12919 1962 12923 1966
rect 12932 1954 12936 1958
rect 12943 1962 12947 1966
rect 12955 1954 12960 1959
rect 12970 1954 12974 1958
rect 12999 1954 13004 1959
rect 13051 1959 13055 1964
rect 13014 1954 13018 1958
rect 9019 1850 9023 1854
rect 9030 1857 9034 1861
rect 9061 1858 9065 1862
rect 8040 1760 8044 1764
rect 8053 1752 8057 1756
rect 8064 1760 8068 1764
rect 8076 1752 8081 1757
rect 8091 1752 8095 1756
rect 8120 1752 8125 1757
rect 8172 1757 8176 1762
rect 8135 1752 8139 1756
rect 8523 1720 8527 1724
rect 8523 1665 8527 1669
rect 8592 1694 8596 1698
rect 8603 1683 8607 1687
rect 8044 1598 8048 1602
rect 8057 1590 8061 1594
rect 8068 1598 8072 1602
rect 8080 1590 8085 1595
rect 8095 1590 8099 1594
rect 8124 1590 8129 1595
rect 8176 1595 8180 1600
rect 8139 1590 8143 1594
rect 9021 1500 9025 1504
rect 9032 1507 9036 1511
rect 12904 1521 12908 1525
rect 9063 1508 9067 1512
rect 12917 1513 12921 1517
rect 12928 1521 12932 1525
rect 12940 1513 12945 1518
rect 12955 1513 12959 1517
rect 12984 1513 12989 1518
rect 13036 1518 13040 1523
rect 12999 1513 13003 1517
rect 12534 1406 12538 1410
rect 8550 1361 8554 1365
rect 8049 1348 8053 1352
rect 8062 1340 8066 1344
rect 8073 1348 8077 1352
rect 8085 1340 8090 1345
rect 8100 1340 8104 1344
rect 8129 1340 8134 1345
rect 8181 1345 8185 1350
rect 8144 1340 8148 1344
rect 12534 1351 12538 1355
rect 8550 1306 8554 1310
rect 8619 1335 8623 1339
rect 12603 1380 12607 1384
rect 12614 1369 12618 1373
rect 8630 1324 8634 1328
rect 9029 1208 9033 1212
rect 9040 1215 9044 1219
rect 9071 1216 9075 1220
rect 8047 1188 8051 1192
rect 8060 1180 8064 1184
rect 8071 1188 8075 1192
rect 8083 1180 8088 1185
rect 8098 1180 8102 1184
rect 8127 1180 8132 1185
rect 8179 1185 8183 1190
rect 8142 1180 8146 1184
rect 8543 1018 8547 1022
rect 8075 953 8079 957
rect 8088 945 8092 949
rect 8099 953 8103 957
rect 8111 945 8116 950
rect 8126 945 8130 949
rect 8155 945 8160 950
rect 8207 950 8211 955
rect 8170 945 8174 949
rect 8543 963 8547 967
rect 8612 992 8616 996
rect 8623 981 8627 985
rect 12474 976 12478 980
rect 12889 968 12893 972
rect 12474 921 12478 925
rect 12543 950 12547 954
rect 12902 960 12906 964
rect 12913 968 12917 972
rect 12925 960 12930 965
rect 12940 960 12944 964
rect 12969 960 12974 965
rect 13021 965 13025 970
rect 12984 960 12988 964
rect 12554 939 12558 943
rect 9017 842 9021 846
rect 9028 849 9032 853
rect 9059 850 9063 854
rect 8084 828 8088 832
rect 8097 820 8101 824
rect 8108 828 8112 832
rect 8120 820 8125 825
rect 8135 820 8139 824
rect 8164 820 8169 825
rect 8216 825 8220 830
rect 8179 820 8183 824
rect 12902 676 12906 680
rect 12915 668 12919 672
rect 12926 676 12930 680
rect 12938 668 12943 673
rect 12953 668 12957 672
rect 12982 668 12987 673
rect 13034 673 13038 678
rect 12997 668 13001 672
rect 12431 440 12435 444
rect 12431 385 12435 389
rect 12500 414 12504 418
rect 12511 403 12515 407
rect 12924 302 12928 306
rect 12937 294 12941 298
rect 12948 302 12952 306
rect 12960 294 12965 299
rect 12975 294 12979 298
rect 13004 294 13009 299
rect 13056 299 13060 304
rect 13019 294 13023 298
<< metal1 >>
rect 7996 2467 8149 2471
rect 8002 2461 8006 2467
rect 8040 2461 8044 2467
rect 8084 2461 8088 2467
rect 8129 2461 8133 2467
rect 8052 2436 8065 2461
rect 8096 2436 8109 2461
rect 7991 2425 7998 2429
rect 8002 2417 8011 2421
rect 8018 2414 8022 2436
rect 8026 2425 8027 2429
rect 8062 2427 8065 2436
rect 8106 2427 8109 2436
rect 8062 2422 8074 2427
rect 8106 2422 8130 2427
rect 8137 2426 8141 2436
rect 8026 2420 8034 2422
rect 8031 2417 8034 2420
rect 8053 2417 8054 2421
rect 8062 2414 8065 2422
rect 8070 2417 8078 2422
rect 8097 2417 8098 2421
rect 8106 2414 8109 2422
rect 8137 2421 8150 2426
rect 8137 2414 8141 2421
rect 8010 2404 8022 2414
rect 8054 2404 8065 2414
rect 8098 2404 8109 2414
rect 7998 2399 8002 2404
rect 8034 2399 8038 2404
rect 8078 2399 8082 2404
rect 8129 2399 8133 2404
rect 7997 2395 8141 2399
rect 7990 2298 8143 2302
rect 7996 2292 8000 2298
rect 8034 2292 8038 2298
rect 8078 2292 8082 2298
rect 8123 2292 8127 2298
rect 8046 2267 8059 2292
rect 8090 2267 8103 2292
rect 7985 2256 7992 2260
rect 7996 2248 8005 2252
rect 8012 2245 8016 2267
rect 8020 2256 8021 2260
rect 8056 2258 8059 2267
rect 8100 2258 8103 2267
rect 8056 2253 8068 2258
rect 8100 2253 8124 2258
rect 8131 2257 8135 2267
rect 8020 2251 8028 2253
rect 8025 2248 8028 2251
rect 8047 2248 8048 2252
rect 8056 2245 8059 2253
rect 8064 2248 8072 2253
rect 8091 2248 8092 2252
rect 8100 2245 8103 2253
rect 8131 2252 8144 2257
rect 8131 2245 8135 2252
rect 12492 2245 12520 2248
rect 8004 2235 8016 2245
rect 8048 2235 8059 2245
rect 8092 2235 8103 2245
rect 12493 2239 12496 2245
rect 12517 2244 12520 2245
rect 12517 2241 12588 2244
rect 7992 2230 7996 2235
rect 8028 2230 8032 2235
rect 8072 2230 8076 2235
rect 8123 2230 8127 2235
rect 7991 2226 8135 2230
rect 12476 2215 12479 2218
rect 12484 2216 12494 2219
rect 12502 2219 12505 2227
rect 12532 2235 12535 2241
rect 12551 2235 12554 2241
rect 12502 2216 12523 2219
rect 12502 2213 12505 2216
rect 12493 2203 12496 2207
rect 12487 2201 12511 2203
rect 12487 2200 12505 2201
rect 12510 2200 12511 2201
rect 12520 2193 12523 2216
rect 12561 2235 12581 2238
rect 12561 2229 12564 2235
rect 12578 2229 12581 2235
rect 12542 2208 12545 2211
rect 12542 2205 12560 2208
rect 12570 2198 12573 2205
rect 12570 2195 12587 2198
rect 12492 2192 12511 2193
rect 12487 2190 12511 2192
rect 12520 2190 12563 2193
rect 12493 2184 12496 2190
rect 12584 2184 12587 2195
rect 12549 2179 12574 2182
rect 12584 2180 12597 2184
rect 12549 2177 12552 2179
rect 12476 2161 12479 2164
rect 12484 2161 12494 2164
rect 12502 2164 12505 2172
rect 12514 2174 12552 2177
rect 12584 2176 12587 2180
rect 12514 2164 12517 2174
rect 12555 2173 12587 2176
rect 12555 2170 12558 2173
rect 12502 2161 12517 2164
rect 12502 2158 12505 2161
rect 12554 2167 12560 2170
rect 12493 2148 12496 2152
rect 12514 2151 12519 2154
rect 12532 2154 12535 2158
rect 12579 2154 12582 2158
rect 12524 2151 12588 2154
rect 12514 2148 12517 2151
rect 12487 2145 12517 2148
rect 12593 2140 12597 2180
rect 7990 2118 8143 2122
rect 7996 2112 8000 2118
rect 8034 2112 8038 2118
rect 8078 2112 8082 2118
rect 8123 2112 8127 2118
rect 8046 2087 8059 2112
rect 8090 2087 8103 2112
rect 8530 2108 8558 2111
rect 8531 2102 8534 2108
rect 8555 2107 8558 2108
rect 8555 2104 8626 2107
rect 7985 2076 7992 2080
rect 7996 2068 8005 2072
rect 8012 2065 8016 2087
rect 8020 2076 8021 2080
rect 8056 2078 8059 2087
rect 8100 2078 8103 2087
rect 8056 2073 8068 2078
rect 8100 2073 8124 2078
rect 8131 2077 8135 2087
rect 8514 2078 8517 2081
rect 8522 2079 8532 2082
rect 8540 2082 8543 2090
rect 8570 2098 8573 2104
rect 8589 2098 8592 2104
rect 8540 2079 8561 2082
rect 8020 2071 8028 2073
rect 8025 2068 8028 2071
rect 8047 2068 8048 2072
rect 8056 2065 8059 2073
rect 8064 2068 8072 2073
rect 8091 2068 8092 2072
rect 8100 2065 8103 2073
rect 8131 2072 8144 2077
rect 8540 2076 8543 2079
rect 8131 2065 8135 2072
rect 8531 2066 8534 2070
rect 8004 2055 8016 2065
rect 8048 2055 8059 2065
rect 8092 2055 8103 2065
rect 8525 2064 8549 2066
rect 8525 2063 8543 2064
rect 8548 2063 8549 2064
rect 8558 2056 8561 2079
rect 8599 2098 8619 2101
rect 8599 2092 8602 2098
rect 8616 2092 8619 2098
rect 8580 2071 8583 2074
rect 8580 2068 8598 2071
rect 8608 2061 8611 2068
rect 13408 2063 13412 2066
rect 8608 2058 8625 2061
rect 13402 2059 13403 2063
rect 13407 2059 13412 2063
rect 8530 2055 8549 2056
rect 7992 2050 7996 2055
rect 8028 2050 8032 2055
rect 8072 2050 8076 2055
rect 8123 2050 8127 2055
rect 8525 2053 8549 2055
rect 8558 2053 8601 2056
rect 7991 2046 8135 2050
rect 8531 2047 8534 2053
rect 8622 2047 8625 2058
rect 13408 2053 13412 2059
rect 8587 2042 8612 2045
rect 8622 2043 8635 2047
rect 8587 2040 8590 2042
rect 8514 2024 8517 2027
rect 8522 2024 8532 2027
rect 8540 2027 8543 2035
rect 8552 2037 8590 2040
rect 8622 2039 8625 2043
rect 8552 2027 8555 2037
rect 8593 2036 8625 2039
rect 8593 2033 8596 2036
rect 8540 2024 8555 2027
rect 8540 2021 8543 2024
rect 8592 2030 8598 2033
rect 8531 2011 8534 2015
rect 8552 2014 8557 2017
rect 8570 2017 8573 2021
rect 8617 2017 8620 2021
rect 8562 2014 8626 2017
rect 8552 2011 8555 2014
rect 8525 2008 8555 2011
rect 8631 2003 8635 2043
rect 10229 2015 10233 2024
rect 10279 2016 10283 2025
rect 10329 2016 10333 2025
rect 10376 2016 10380 2025
rect 13416 2023 13420 2033
rect 13416 2019 13425 2023
rect 10223 2010 10224 2015
rect 10228 2010 10247 2015
rect 10273 2011 10274 2016
rect 10278 2011 10297 2016
rect 10323 2011 10324 2016
rect 10328 2011 10347 2016
rect 10370 2011 10371 2016
rect 10375 2011 10394 2016
rect 13416 2015 13420 2019
rect 10229 2004 10233 2010
rect 10279 2005 10283 2011
rect 10329 2005 10333 2011
rect 10376 2005 10380 2011
rect 12917 2004 13070 2008
rect 12923 1998 12927 2004
rect 12961 1998 12965 2004
rect 13005 1998 13009 2004
rect 13050 1998 13054 2004
rect 12973 1973 12986 1998
rect 13017 1973 13030 1998
rect 13408 1995 13412 2005
rect 12912 1962 12919 1966
rect 10237 1940 10241 1954
rect 10287 1941 10291 1955
rect 10337 1941 10341 1955
rect 10384 1941 10388 1955
rect 12923 1954 12932 1958
rect 12939 1951 12943 1973
rect 12947 1962 12948 1966
rect 12983 1964 12986 1973
rect 13027 1964 13030 1973
rect 12983 1959 12995 1964
rect 13027 1959 13051 1964
rect 13058 1963 13062 1973
rect 12947 1957 12955 1959
rect 12952 1954 12955 1957
rect 12974 1954 12975 1958
rect 12983 1951 12986 1959
rect 12991 1954 12999 1959
rect 13018 1954 13019 1958
rect 13027 1951 13030 1959
rect 13058 1958 13071 1963
rect 13058 1951 13062 1958
rect 12931 1941 12943 1951
rect 12975 1941 12986 1951
rect 13019 1941 13030 1951
rect 12919 1936 12923 1941
rect 12955 1936 12959 1941
rect 12999 1936 13003 1941
rect 13050 1936 13054 1941
rect 12918 1932 13062 1936
rect 9018 1907 9041 1911
rect 9022 1905 9041 1907
rect 9018 1896 9022 1901
rect 9037 1896 9041 1905
rect 9054 1900 9078 1901
rect 9054 1896 9070 1900
rect 9074 1896 9078 1900
rect 9054 1894 9078 1896
rect 9060 1889 9064 1894
rect 9029 1868 9033 1876
rect 9029 1864 9041 1868
rect 9037 1862 9041 1864
rect 9068 1862 9072 1869
rect 9012 1857 9030 1861
rect 9037 1858 9061 1862
rect 9068 1858 9078 1862
rect 9012 1850 9019 1854
rect 9037 1847 9041 1858
rect 9068 1855 9072 1858
rect 9060 1841 9064 1845
rect 9054 1840 9079 1841
rect 9054 1836 9074 1840
rect 9054 1835 9079 1836
rect 9018 1823 9022 1827
rect 9018 1819 9034 1823
rect 8038 1802 8191 1806
rect 8044 1796 8048 1802
rect 8082 1796 8086 1802
rect 8126 1796 8130 1802
rect 8171 1796 8175 1802
rect 8094 1771 8107 1796
rect 8138 1771 8151 1796
rect 10698 1786 10718 1790
rect 10729 1786 10760 1790
rect 10772 1786 10800 1790
rect 10810 1786 10831 1790
rect 10847 1788 10877 1792
rect 10698 1783 10702 1786
rect 10736 1783 10740 1786
rect 10780 1783 10784 1786
rect 10818 1783 10822 1786
rect 10864 1785 10868 1788
rect 10692 1779 10693 1783
rect 10697 1779 10702 1783
rect 10730 1779 10731 1783
rect 10735 1779 10740 1783
rect 10774 1779 10775 1783
rect 10779 1779 10784 1783
rect 10812 1779 10813 1783
rect 10817 1779 10822 1783
rect 10858 1781 10859 1785
rect 10863 1781 10868 1785
rect 8033 1760 8040 1764
rect 8044 1752 8053 1756
rect 8060 1749 8064 1771
rect 8068 1760 8069 1764
rect 8104 1762 8107 1771
rect 8148 1762 8151 1771
rect 8104 1757 8116 1762
rect 8148 1757 8172 1762
rect 8179 1761 8183 1771
rect 10165 1768 10169 1776
rect 10193 1768 10197 1776
rect 10220 1768 10224 1776
rect 10259 1768 10263 1776
rect 10287 1768 10291 1776
rect 10314 1768 10318 1776
rect 10354 1769 10358 1777
rect 10382 1769 10386 1777
rect 10409 1769 10413 1777
rect 10445 1769 10449 1777
rect 10698 1773 10702 1779
rect 10736 1773 10740 1779
rect 10780 1773 10784 1779
rect 10818 1773 10822 1779
rect 10864 1775 10868 1781
rect 8068 1755 8076 1757
rect 8073 1752 8076 1755
rect 8095 1752 8096 1756
rect 8104 1749 8107 1757
rect 8112 1752 8120 1757
rect 8139 1752 8140 1756
rect 8148 1749 8151 1757
rect 8179 1756 8192 1761
rect 8179 1749 8183 1756
rect 8521 1749 8549 1752
rect 8052 1739 8064 1749
rect 8096 1739 8107 1749
rect 8140 1739 8151 1749
rect 8522 1743 8525 1749
rect 8546 1748 8549 1749
rect 8546 1745 8617 1748
rect 8040 1734 8044 1739
rect 8076 1734 8080 1739
rect 8120 1734 8124 1739
rect 8171 1734 8175 1739
rect 8039 1730 8183 1734
rect 8505 1719 8508 1722
rect 8513 1720 8523 1723
rect 8531 1723 8534 1731
rect 8561 1739 8564 1745
rect 8580 1739 8583 1745
rect 8531 1720 8552 1723
rect 8531 1717 8534 1720
rect 8522 1707 8525 1711
rect 8516 1705 8540 1707
rect 8516 1704 8534 1705
rect 8539 1704 8540 1705
rect 8549 1697 8552 1720
rect 8590 1739 8610 1742
rect 8590 1733 8593 1739
rect 8607 1733 8610 1739
rect 8571 1712 8574 1715
rect 8571 1709 8589 1712
rect 8599 1702 8602 1709
rect 8599 1699 8616 1702
rect 8521 1696 8540 1697
rect 8516 1694 8540 1696
rect 8549 1694 8592 1697
rect 8522 1688 8525 1694
rect 8613 1688 8616 1699
rect 8578 1683 8603 1686
rect 8613 1684 8626 1688
rect 8578 1681 8581 1683
rect 8505 1665 8508 1668
rect 8513 1665 8523 1668
rect 8531 1668 8534 1676
rect 8543 1678 8581 1681
rect 8613 1680 8616 1684
rect 8543 1668 8546 1678
rect 8584 1677 8616 1680
rect 8584 1674 8587 1677
rect 8531 1665 8546 1668
rect 8531 1662 8534 1665
rect 8583 1671 8589 1674
rect 8522 1652 8525 1656
rect 8543 1655 8548 1658
rect 8561 1658 8564 1662
rect 8608 1658 8611 1662
rect 8553 1655 8617 1658
rect 8543 1652 8546 1655
rect 8516 1649 8546 1652
rect 8622 1644 8626 1684
rect 10706 1715 10710 1733
rect 10744 1715 10748 1733
rect 10788 1715 10792 1733
rect 10826 1715 10830 1733
rect 10872 1717 10876 1735
rect 10698 1686 10702 1695
rect 10736 1686 10740 1695
rect 10780 1686 10784 1695
rect 10818 1686 10822 1695
rect 10864 1688 10868 1697
rect 10698 1682 10718 1686
rect 10729 1682 10760 1686
rect 10772 1682 10800 1686
rect 10810 1682 10827 1686
rect 10847 1684 10873 1688
rect 10173 1662 10177 1668
rect 10201 1662 10205 1668
rect 10228 1662 10232 1668
rect 10267 1662 10271 1668
rect 10295 1662 10299 1668
rect 10322 1662 10326 1668
rect 10362 1663 10366 1669
rect 10390 1663 10394 1669
rect 10417 1663 10421 1669
rect 10453 1663 10457 1669
rect 8042 1640 8195 1644
rect 13436 1642 13440 1645
rect 8048 1634 8052 1640
rect 8086 1634 8090 1640
rect 8130 1634 8134 1640
rect 8175 1634 8179 1640
rect 13430 1638 13431 1642
rect 13435 1638 13440 1642
rect 8098 1609 8111 1634
rect 8142 1609 8155 1634
rect 13436 1632 13440 1638
rect 8037 1598 8044 1602
rect 8048 1590 8057 1594
rect 8064 1587 8068 1609
rect 8072 1598 8073 1602
rect 8108 1600 8111 1609
rect 8152 1600 8155 1609
rect 8108 1595 8120 1600
rect 8152 1595 8176 1600
rect 8183 1599 8187 1609
rect 13444 1602 13448 1612
rect 8072 1593 8080 1595
rect 8077 1590 8080 1593
rect 8099 1590 8100 1594
rect 8108 1587 8111 1595
rect 8116 1590 8124 1595
rect 8143 1590 8144 1594
rect 8152 1587 8155 1595
rect 8183 1594 8196 1599
rect 13444 1598 13453 1602
rect 13444 1594 13448 1598
rect 8183 1587 8187 1594
rect 8056 1577 8068 1587
rect 8100 1577 8111 1587
rect 8144 1577 8155 1587
rect 8044 1572 8048 1577
rect 8080 1572 8084 1577
rect 8124 1572 8128 1577
rect 8175 1572 8179 1577
rect 13436 1574 13440 1584
rect 8043 1568 8187 1572
rect 12902 1563 13055 1567
rect 9020 1557 9043 1561
rect 9024 1555 9043 1557
rect 9020 1546 9024 1551
rect 9039 1546 9043 1555
rect 12908 1557 12912 1563
rect 12946 1557 12950 1563
rect 12990 1557 12994 1563
rect 13035 1557 13039 1563
rect 9056 1550 9080 1551
rect 9056 1546 9072 1550
rect 9076 1546 9080 1550
rect 9056 1544 9080 1546
rect 9062 1539 9066 1544
rect 9031 1518 9035 1526
rect 12958 1532 12971 1557
rect 13002 1532 13015 1557
rect 12897 1521 12904 1525
rect 9031 1514 9043 1518
rect 9039 1512 9043 1514
rect 9070 1512 9074 1519
rect 12908 1513 12917 1517
rect 9014 1507 9032 1511
rect 9039 1508 9063 1512
rect 9070 1508 9080 1512
rect 12924 1510 12928 1532
rect 12932 1521 12933 1525
rect 12968 1523 12971 1532
rect 13012 1523 13015 1532
rect 12968 1518 12980 1523
rect 13012 1518 13036 1523
rect 13043 1522 13047 1532
rect 12932 1516 12940 1518
rect 12937 1513 12940 1516
rect 12959 1513 12960 1517
rect 12968 1510 12971 1518
rect 12976 1513 12984 1518
rect 13003 1513 13004 1517
rect 13012 1510 13015 1518
rect 13043 1517 13056 1522
rect 13043 1510 13047 1517
rect 9014 1500 9021 1504
rect 9039 1497 9043 1508
rect 9070 1505 9074 1508
rect 12916 1500 12928 1510
rect 12960 1500 12971 1510
rect 13004 1500 13015 1510
rect 12904 1495 12908 1500
rect 12940 1495 12944 1500
rect 12984 1495 12988 1500
rect 13035 1495 13039 1500
rect 9062 1491 9066 1495
rect 12903 1491 13047 1495
rect 9056 1490 9081 1491
rect 9056 1486 9076 1490
rect 9056 1485 9081 1486
rect 9020 1473 9024 1477
rect 9020 1469 9036 1473
rect 12532 1435 12560 1438
rect 12533 1429 12536 1435
rect 12557 1434 12560 1435
rect 12557 1431 12628 1434
rect 12516 1405 12519 1408
rect 12524 1406 12534 1409
rect 12542 1409 12545 1417
rect 12572 1425 12575 1431
rect 12591 1425 12594 1431
rect 12542 1406 12563 1409
rect 12542 1403 12545 1406
rect 8047 1390 8200 1394
rect 12533 1393 12536 1397
rect 8548 1390 8576 1393
rect 12527 1391 12551 1393
rect 12527 1390 12545 1391
rect 8053 1384 8057 1390
rect 8091 1384 8095 1390
rect 8135 1384 8139 1390
rect 8180 1384 8184 1390
rect 8549 1384 8552 1390
rect 8573 1389 8576 1390
rect 8573 1386 8644 1389
rect 8103 1359 8116 1384
rect 8147 1359 8160 1384
rect 8532 1360 8535 1363
rect 8540 1361 8550 1364
rect 8558 1364 8561 1372
rect 8588 1380 8591 1386
rect 8607 1380 8610 1386
rect 8558 1361 8579 1364
rect 8042 1348 8049 1352
rect 8053 1340 8062 1344
rect 8069 1337 8073 1359
rect 8077 1348 8078 1352
rect 8113 1350 8116 1359
rect 8157 1350 8160 1359
rect 8113 1345 8125 1350
rect 8157 1345 8181 1350
rect 8188 1349 8192 1359
rect 8558 1358 8561 1361
rect 8077 1343 8085 1345
rect 8082 1340 8085 1343
rect 8104 1340 8105 1344
rect 8113 1337 8116 1345
rect 8121 1340 8129 1345
rect 8148 1340 8149 1344
rect 8157 1337 8160 1345
rect 8188 1344 8201 1349
rect 8549 1348 8552 1352
rect 8543 1346 8567 1348
rect 8543 1345 8561 1346
rect 8188 1337 8192 1344
rect 8061 1327 8073 1337
rect 8105 1327 8116 1337
rect 8149 1327 8160 1337
rect 8566 1345 8567 1346
rect 8576 1338 8579 1361
rect 8617 1380 8637 1383
rect 12550 1390 12551 1391
rect 12560 1383 12563 1406
rect 12601 1425 12621 1428
rect 12601 1419 12604 1425
rect 12618 1419 12621 1425
rect 12582 1398 12585 1401
rect 12582 1395 12600 1398
rect 12610 1388 12613 1395
rect 12610 1385 12627 1388
rect 12532 1382 12551 1383
rect 12527 1380 12551 1382
rect 12560 1380 12603 1383
rect 8617 1374 8620 1380
rect 8634 1374 8637 1380
rect 12533 1374 12536 1380
rect 12624 1374 12627 1385
rect 8598 1353 8601 1356
rect 8598 1350 8616 1353
rect 12589 1369 12614 1372
rect 12624 1370 12637 1374
rect 12589 1367 12592 1369
rect 12516 1351 12519 1354
rect 12524 1351 12534 1354
rect 12542 1354 12545 1362
rect 12554 1364 12592 1367
rect 12624 1366 12627 1370
rect 12554 1354 12557 1364
rect 12595 1363 12627 1366
rect 12595 1360 12598 1363
rect 12542 1351 12557 1354
rect 8626 1343 8629 1350
rect 12542 1348 12545 1351
rect 8626 1340 8643 1343
rect 8548 1337 8567 1338
rect 8543 1335 8567 1337
rect 8576 1335 8619 1338
rect 8549 1329 8552 1335
rect 8640 1329 8643 1340
rect 12594 1357 12600 1360
rect 12533 1338 12536 1342
rect 12554 1341 12559 1344
rect 12572 1344 12575 1348
rect 12619 1344 12622 1348
rect 12564 1341 12628 1344
rect 12554 1338 12557 1341
rect 12527 1335 12557 1338
rect 12633 1330 12637 1370
rect 8049 1322 8053 1327
rect 8085 1322 8089 1327
rect 8129 1322 8133 1327
rect 8180 1322 8184 1327
rect 8048 1318 8192 1322
rect 8605 1324 8630 1327
rect 8640 1325 8653 1329
rect 8605 1322 8608 1324
rect 8532 1306 8535 1309
rect 8540 1306 8550 1309
rect 8558 1309 8561 1317
rect 8570 1319 8608 1322
rect 8640 1321 8643 1325
rect 8570 1309 8573 1319
rect 8611 1318 8643 1321
rect 8611 1315 8614 1318
rect 8558 1306 8573 1309
rect 8558 1303 8561 1306
rect 8610 1312 8616 1315
rect 8549 1293 8552 1297
rect 8570 1296 8575 1299
rect 8588 1299 8591 1303
rect 8635 1299 8638 1303
rect 8580 1296 8644 1299
rect 8570 1293 8573 1296
rect 8543 1290 8573 1293
rect 8649 1285 8653 1325
rect 9028 1265 9051 1269
rect 9032 1263 9051 1265
rect 9028 1254 9032 1259
rect 9047 1254 9051 1263
rect 9064 1258 9088 1259
rect 9064 1254 9080 1258
rect 9084 1254 9088 1258
rect 9064 1252 9088 1254
rect 9070 1247 9074 1252
rect 8045 1230 8198 1234
rect 8051 1224 8055 1230
rect 8089 1224 8093 1230
rect 8133 1224 8137 1230
rect 8178 1224 8182 1230
rect 9039 1226 9043 1234
rect 8101 1199 8114 1224
rect 8145 1199 8158 1224
rect 9039 1222 9051 1226
rect 9047 1220 9051 1222
rect 9078 1220 9082 1227
rect 9022 1215 9040 1219
rect 9047 1216 9071 1220
rect 9078 1216 9088 1220
rect 9022 1208 9029 1212
rect 9047 1205 9051 1216
rect 9078 1213 9082 1216
rect 8040 1188 8047 1192
rect 8051 1180 8060 1184
rect 8067 1177 8071 1199
rect 8075 1188 8076 1192
rect 8111 1190 8114 1199
rect 8155 1190 8158 1199
rect 8111 1185 8123 1190
rect 8155 1185 8179 1190
rect 8186 1189 8190 1199
rect 8075 1183 8083 1185
rect 8080 1180 8083 1183
rect 8102 1180 8103 1184
rect 8111 1177 8114 1185
rect 8119 1180 8127 1185
rect 8146 1180 8147 1184
rect 8155 1177 8158 1185
rect 8186 1184 8199 1189
rect 9070 1199 9074 1203
rect 9064 1198 9089 1199
rect 9064 1194 9084 1198
rect 9064 1193 9089 1194
rect 8186 1177 8190 1184
rect 9028 1181 9032 1185
rect 9028 1177 9044 1181
rect 8059 1167 8071 1177
rect 8103 1167 8114 1177
rect 8147 1167 8158 1177
rect 8047 1162 8051 1167
rect 8083 1162 8087 1167
rect 8127 1162 8131 1167
rect 8178 1162 8182 1167
rect 8046 1158 8190 1162
rect 13487 1088 13491 1091
rect 13481 1084 13482 1088
rect 13486 1084 13491 1088
rect 13487 1078 13491 1084
rect 8541 1047 8569 1050
rect 13495 1048 13499 1058
rect 8542 1041 8545 1047
rect 8566 1046 8569 1047
rect 8566 1043 8637 1046
rect 13495 1044 13504 1048
rect 8525 1017 8528 1020
rect 8533 1018 8543 1021
rect 8551 1021 8554 1029
rect 8581 1037 8584 1043
rect 8600 1037 8603 1043
rect 13495 1040 13499 1044
rect 8551 1018 8572 1021
rect 8551 1015 8554 1018
rect 8542 1005 8545 1009
rect 8536 1003 8560 1005
rect 8536 1002 8554 1003
rect 8073 995 8226 999
rect 8079 989 8083 995
rect 8117 989 8121 995
rect 8161 989 8165 995
rect 8206 989 8210 995
rect 8559 1002 8560 1003
rect 8569 995 8572 1018
rect 8610 1037 8630 1040
rect 8610 1031 8613 1037
rect 8627 1031 8630 1037
rect 8591 1010 8594 1013
rect 8591 1007 8609 1010
rect 13487 1020 13491 1030
rect 12887 1010 13040 1014
rect 8619 1000 8622 1007
rect 12472 1005 12500 1008
rect 8619 997 8636 1000
rect 8541 994 8560 995
rect 8536 992 8560 994
rect 8569 992 8612 995
rect 8129 964 8142 989
rect 8173 964 8186 989
rect 8542 986 8545 992
rect 8633 986 8636 997
rect 12473 999 12476 1005
rect 12497 1004 12500 1005
rect 12893 1004 12897 1010
rect 12931 1004 12935 1010
rect 12975 1004 12979 1010
rect 13020 1004 13024 1010
rect 12497 1001 12568 1004
rect 8598 981 8623 984
rect 8633 982 8646 986
rect 8598 979 8601 981
rect 8068 953 8075 957
rect 8079 945 8088 949
rect 8095 942 8099 964
rect 8103 953 8104 957
rect 8139 955 8142 964
rect 8183 955 8186 964
rect 8139 950 8151 955
rect 8183 950 8207 955
rect 8214 954 8218 964
rect 8525 963 8528 966
rect 8533 963 8543 966
rect 8551 966 8554 974
rect 8563 976 8601 979
rect 8633 978 8636 982
rect 8563 966 8566 976
rect 8604 975 8636 978
rect 8604 972 8607 975
rect 8551 963 8566 966
rect 8551 960 8554 963
rect 8603 969 8609 972
rect 8103 948 8111 950
rect 8108 945 8111 948
rect 8130 945 8131 949
rect 8139 942 8142 950
rect 8147 945 8155 950
rect 8174 945 8175 949
rect 8183 942 8186 950
rect 8214 949 8227 954
rect 8542 950 8545 954
rect 8563 953 8568 956
rect 8581 956 8584 960
rect 8628 956 8631 960
rect 8573 953 8637 956
rect 8563 950 8566 953
rect 8214 942 8218 949
rect 8536 947 8566 950
rect 8642 942 8646 982
rect 12456 975 12459 978
rect 12464 976 12474 979
rect 12482 979 12485 987
rect 12512 995 12515 1001
rect 12531 995 12534 1001
rect 12482 976 12503 979
rect 12482 973 12485 976
rect 12473 963 12476 967
rect 12467 961 12491 963
rect 12467 960 12485 961
rect 12490 960 12491 961
rect 12500 953 12503 976
rect 12541 995 12561 998
rect 12541 989 12544 995
rect 12558 989 12561 995
rect 12522 968 12525 971
rect 12522 965 12540 968
rect 12943 979 12956 1004
rect 12987 979 13000 1004
rect 12882 968 12889 972
rect 12550 958 12553 965
rect 12893 960 12902 964
rect 12550 955 12567 958
rect 12909 957 12913 979
rect 12917 968 12918 972
rect 12953 970 12956 979
rect 12997 970 13000 979
rect 12953 965 12965 970
rect 12997 965 13021 970
rect 13028 969 13032 979
rect 12917 963 12925 965
rect 12922 960 12925 963
rect 12944 960 12945 964
rect 12953 957 12956 965
rect 12961 960 12969 965
rect 12988 960 12989 964
rect 12997 957 13000 965
rect 13028 964 13041 969
rect 13028 957 13032 964
rect 12472 952 12491 953
rect 12467 950 12491 952
rect 12500 950 12543 953
rect 12473 944 12476 950
rect 12564 944 12567 955
rect 12901 947 12913 957
rect 12945 947 12956 957
rect 12989 947 13000 957
rect 8087 932 8099 942
rect 8131 932 8142 942
rect 8175 932 8186 942
rect 12529 939 12554 942
rect 12564 940 12577 944
rect 12889 942 12893 947
rect 12925 942 12929 947
rect 12969 942 12973 947
rect 13020 942 13024 947
rect 12529 937 12532 939
rect 8075 927 8079 932
rect 8111 927 8115 932
rect 8155 927 8159 932
rect 8206 927 8210 932
rect 8074 923 8218 927
rect 12456 921 12459 924
rect 12464 921 12474 924
rect 12482 924 12485 932
rect 12494 934 12532 937
rect 12564 936 12567 940
rect 12494 924 12497 934
rect 12535 933 12567 936
rect 12535 930 12538 933
rect 12482 921 12497 924
rect 12482 918 12485 921
rect 12534 927 12540 930
rect 12473 908 12476 912
rect 12494 911 12499 914
rect 12512 914 12515 918
rect 12559 914 12562 918
rect 12504 911 12568 914
rect 12494 908 12497 911
rect 12467 905 12497 908
rect 9016 899 9039 903
rect 12573 900 12577 940
rect 12888 938 13032 942
rect 9020 897 9039 899
rect 9016 888 9020 893
rect 9035 888 9039 897
rect 8082 870 8235 874
rect 8088 864 8092 870
rect 8126 864 8130 870
rect 8170 864 8174 870
rect 8215 864 8219 870
rect 9052 892 9076 893
rect 9052 888 9068 892
rect 9072 888 9076 892
rect 9052 886 9076 888
rect 9058 881 9062 886
rect 8138 839 8151 864
rect 8182 839 8195 864
rect 9027 860 9031 868
rect 9027 856 9039 860
rect 9035 854 9039 856
rect 9066 854 9070 861
rect 9010 849 9028 853
rect 9035 850 9059 854
rect 9066 850 9076 854
rect 9010 842 9017 846
rect 9035 839 9039 850
rect 9066 847 9070 850
rect 8077 828 8084 832
rect 8088 820 8097 824
rect 8104 817 8108 839
rect 8112 828 8113 832
rect 8148 830 8151 839
rect 8192 830 8195 839
rect 8148 825 8160 830
rect 8192 825 8216 830
rect 8223 829 8227 839
rect 8112 823 8120 825
rect 8117 820 8120 823
rect 8139 820 8140 824
rect 8148 817 8151 825
rect 8156 820 8164 825
rect 8183 820 8184 824
rect 8192 817 8195 825
rect 8223 824 8236 829
rect 8223 817 8227 824
rect 8096 807 8108 817
rect 8140 807 8151 817
rect 8184 807 8195 817
rect 9058 833 9062 837
rect 9052 832 9077 833
rect 9052 828 9072 832
rect 9052 827 9077 828
rect 9016 815 9020 819
rect 9016 811 9032 815
rect 8084 802 8088 807
rect 8120 802 8124 807
rect 8164 802 8168 807
rect 8215 802 8219 807
rect 8083 798 8227 802
rect 13472 739 13476 742
rect 13466 735 13467 739
rect 13471 735 13476 739
rect 13472 729 13476 735
rect 12900 718 13053 722
rect 12906 712 12910 718
rect 12944 712 12948 718
rect 12988 712 12992 718
rect 13033 712 13037 718
rect 12956 687 12969 712
rect 13000 687 13013 712
rect 13480 699 13484 709
rect 13480 695 13489 699
rect 13480 691 13484 695
rect 12895 676 12902 680
rect 12906 668 12915 672
rect 12922 665 12926 687
rect 12930 676 12931 680
rect 12966 678 12969 687
rect 13010 678 13013 687
rect 12966 673 12978 678
rect 13010 673 13034 678
rect 13041 677 13045 687
rect 12930 671 12938 673
rect 12935 668 12938 671
rect 12957 668 12958 672
rect 12966 665 12969 673
rect 12974 668 12982 673
rect 13001 668 13002 672
rect 13010 665 13013 673
rect 13041 672 13054 677
rect 13041 665 13045 672
rect 13472 671 13476 681
rect 12914 655 12926 665
rect 12958 655 12969 665
rect 13002 655 13013 665
rect 12902 650 12906 655
rect 12938 650 12942 655
rect 12982 650 12986 655
rect 13033 650 13037 655
rect 12901 646 13045 650
rect 12429 469 12457 472
rect 12430 463 12433 469
rect 12454 468 12457 469
rect 12454 465 12525 468
rect 12413 439 12416 442
rect 12421 440 12431 443
rect 12439 443 12442 451
rect 12469 459 12472 465
rect 12488 459 12491 465
rect 12439 440 12460 443
rect 12439 437 12442 440
rect 12430 427 12433 431
rect 12424 425 12448 427
rect 12424 424 12442 425
rect 12447 424 12448 425
rect 12457 417 12460 440
rect 12498 459 12518 462
rect 12498 453 12501 459
rect 12515 453 12518 459
rect 12479 432 12482 435
rect 12479 429 12497 432
rect 12507 422 12510 429
rect 12507 419 12524 422
rect 12429 416 12448 417
rect 12424 414 12448 416
rect 12457 414 12500 417
rect 12430 408 12433 414
rect 12521 408 12524 419
rect 12486 403 12511 406
rect 12521 404 12534 408
rect 12486 401 12489 403
rect 12413 385 12416 388
rect 12421 385 12431 388
rect 12439 388 12442 396
rect 12451 398 12489 401
rect 12521 400 12524 404
rect 12451 388 12454 398
rect 12492 397 12524 400
rect 12492 394 12495 397
rect 12439 385 12454 388
rect 12439 382 12442 385
rect 12491 391 12497 394
rect 12430 372 12433 376
rect 12451 375 12456 378
rect 12469 378 12472 382
rect 12516 378 12519 382
rect 12461 375 12525 378
rect 12451 372 12454 375
rect 12424 369 12454 372
rect 12530 364 12534 404
rect 13525 354 13529 357
rect 13519 350 13520 354
rect 13524 350 13529 354
rect 12922 344 13075 348
rect 13525 344 13529 350
rect 12928 338 12932 344
rect 12966 338 12970 344
rect 13010 338 13014 344
rect 13055 338 13059 344
rect 12978 313 12991 338
rect 13022 313 13035 338
rect 13533 314 13537 324
rect 12917 302 12924 306
rect 12928 294 12937 298
rect 12944 291 12948 313
rect 12952 302 12953 306
rect 12988 304 12991 313
rect 13032 304 13035 313
rect 12988 299 13000 304
rect 13032 299 13056 304
rect 13063 303 13067 313
rect 13533 310 13542 314
rect 13533 306 13537 310
rect 12952 297 12960 299
rect 12957 294 12960 297
rect 12979 294 12980 298
rect 12988 291 12991 299
rect 12996 294 13004 299
rect 13023 294 13024 298
rect 13032 291 13035 299
rect 13063 298 13076 303
rect 13063 291 13067 298
rect 12936 281 12948 291
rect 12980 281 12991 291
rect 13024 281 13035 291
rect 13525 286 13529 296
rect 12924 276 12928 281
rect 12960 276 12964 281
rect 13004 276 13008 281
rect 13055 276 13059 281
rect 12923 272 13067 276
<< m2contact >>
rect 7997 2417 8002 2422
rect 8027 2425 8032 2430
rect 8026 2415 8031 2420
rect 8054 2417 8059 2422
rect 8098 2417 8103 2422
rect 7991 2248 7996 2253
rect 8021 2256 8026 2261
rect 8020 2246 8025 2251
rect 8048 2248 8053 2253
rect 8092 2248 8097 2253
rect 12479 2214 12484 2219
rect 12479 2160 12484 2165
rect 7991 2068 7996 2073
rect 8021 2076 8026 2081
rect 8517 2077 8522 2082
rect 8020 2066 8025 2071
rect 8048 2068 8053 2073
rect 8092 2068 8097 2073
rect 8517 2023 8522 2028
rect 12918 1954 12923 1959
rect 12948 1962 12953 1967
rect 12947 1952 12952 1957
rect 12975 1954 12980 1959
rect 13019 1954 13024 1959
rect 8039 1752 8044 1757
rect 8069 1760 8074 1765
rect 8068 1750 8073 1755
rect 8096 1752 8101 1757
rect 8140 1752 8145 1757
rect 8508 1718 8513 1723
rect 8508 1664 8513 1669
rect 8043 1590 8048 1595
rect 8073 1598 8078 1603
rect 8072 1588 8077 1593
rect 8100 1590 8105 1595
rect 8144 1590 8149 1595
rect 12903 1513 12908 1518
rect 12933 1521 12938 1526
rect 12932 1511 12937 1516
rect 12960 1513 12965 1518
rect 13004 1513 13009 1518
rect 12519 1404 12524 1409
rect 8535 1359 8540 1364
rect 8048 1340 8053 1345
rect 8078 1348 8083 1353
rect 8077 1338 8082 1343
rect 8105 1340 8110 1345
rect 8149 1340 8154 1345
rect 12519 1350 12524 1355
rect 8535 1305 8540 1310
rect 8046 1180 8051 1185
rect 8076 1188 8081 1193
rect 8075 1178 8080 1183
rect 8103 1180 8108 1185
rect 8147 1180 8152 1185
rect 8528 1016 8533 1021
rect 8074 945 8079 950
rect 8104 953 8109 958
rect 8528 962 8533 967
rect 8103 943 8108 948
rect 8131 945 8136 950
rect 8175 945 8180 950
rect 12459 974 12464 979
rect 12888 960 12893 965
rect 12918 968 12923 973
rect 12917 958 12922 963
rect 12945 960 12950 965
rect 12989 960 12994 965
rect 12459 920 12464 925
rect 8083 820 8088 825
rect 8113 828 8118 833
rect 8112 818 8117 823
rect 8140 820 8145 825
rect 8184 820 8189 825
rect 12901 668 12906 673
rect 12931 676 12936 681
rect 12930 666 12935 671
rect 12958 668 12963 673
rect 13002 668 13007 673
rect 12416 438 12421 443
rect 12416 384 12421 389
rect 12923 294 12928 299
rect 12953 302 12958 307
rect 12952 292 12957 297
rect 12980 294 12985 299
rect 13024 294 13029 299
<< pm12contact >>
rect 12535 2197 12540 2202
rect 12544 2196 12549 2201
rect 8573 2060 8578 2065
rect 8582 2059 8587 2064
rect 13408 2018 13413 2023
rect 10228 1931 10234 1937
rect 10278 1932 10284 1938
rect 10328 1932 10334 1938
rect 10375 1932 10381 1938
rect 8564 1701 8569 1706
rect 8573 1700 8578 1705
rect 10698 1718 10703 1723
rect 10736 1718 10741 1723
rect 10780 1718 10785 1723
rect 10818 1718 10823 1723
rect 10864 1720 10869 1725
rect 10165 1656 10170 1661
rect 10193 1656 10198 1661
rect 10220 1656 10225 1661
rect 10259 1656 10264 1661
rect 10287 1656 10292 1661
rect 10314 1656 10319 1661
rect 10354 1657 10359 1662
rect 10382 1657 10387 1662
rect 10409 1657 10414 1662
rect 10445 1657 10450 1662
rect 13436 1597 13441 1602
rect 12575 1387 12580 1392
rect 12584 1386 12589 1391
rect 8591 1342 8596 1347
rect 8600 1341 8605 1346
rect 13487 1043 13492 1048
rect 8584 999 8589 1004
rect 8593 998 8598 1003
rect 12515 957 12520 962
rect 12524 956 12529 961
rect 13472 694 13477 699
rect 12472 421 12477 426
rect 12481 420 12486 425
rect 13525 309 13530 314
<< metal2 >>
rect 8027 2475 8058 2478
rect 8027 2430 8031 2475
rect 8054 2422 8058 2475
rect 7976 2417 7997 2421
rect 7988 2393 7994 2417
rect 8027 2393 8031 2415
rect 8098 2393 8103 2417
rect 7988 2390 8107 2393
rect 8021 2306 8052 2309
rect 8021 2261 8025 2306
rect 8048 2253 8052 2306
rect 7970 2248 7991 2252
rect 7982 2224 7988 2248
rect 8021 2224 8025 2246
rect 8092 2224 8097 2248
rect 7982 2221 8101 2224
rect 12480 2208 12483 2214
rect 12480 2205 12517 2208
rect 12514 2202 12517 2205
rect 12514 2199 12535 2202
rect 12544 2186 12547 2196
rect 12481 2183 12547 2186
rect 12481 2165 12484 2183
rect 8021 2126 8052 2129
rect 8021 2081 8025 2126
rect 8048 2073 8052 2126
rect 7970 2068 7991 2072
rect 7982 2044 7988 2068
rect 8518 2071 8521 2077
rect 8518 2068 8555 2071
rect 8021 2044 8025 2066
rect 8092 2044 8097 2068
rect 8552 2065 8555 2068
rect 8552 2062 8573 2065
rect 8582 2049 8585 2059
rect 8519 2046 8585 2049
rect 7982 2041 8101 2044
rect 8519 2028 8522 2046
rect 13399 2018 13408 2023
rect 12948 2012 12979 2015
rect 12948 1967 12952 2012
rect 12975 1959 12979 2012
rect 12897 1954 12918 1958
rect 10218 1931 10228 1937
rect 10268 1932 10278 1938
rect 10318 1932 10328 1938
rect 10365 1932 10375 1938
rect 12909 1930 12915 1954
rect 12948 1930 12952 1952
rect 13019 1930 13024 1954
rect 12909 1927 13028 1930
rect 8069 1810 8100 1813
rect 8069 1765 8073 1810
rect 8096 1757 8100 1810
rect 8018 1752 8039 1756
rect 8030 1728 8036 1752
rect 8069 1728 8073 1750
rect 8140 1728 8145 1752
rect 8030 1725 8149 1728
rect 10695 1718 10698 1723
rect 10733 1718 10736 1723
rect 10777 1718 10780 1723
rect 10815 1718 10818 1723
rect 10861 1720 10864 1725
rect 8509 1712 8512 1718
rect 8509 1709 8546 1712
rect 8543 1706 8546 1709
rect 8543 1703 8564 1706
rect 8573 1690 8576 1700
rect 8510 1687 8576 1690
rect 8510 1669 8513 1687
rect 10161 1656 10165 1661
rect 10189 1656 10193 1661
rect 10216 1656 10220 1661
rect 10255 1656 10259 1661
rect 10283 1656 10287 1661
rect 10310 1656 10314 1661
rect 10350 1657 10354 1662
rect 10378 1657 10382 1662
rect 10405 1657 10409 1662
rect 10441 1657 10445 1662
rect 8073 1648 8104 1651
rect 8073 1603 8077 1648
rect 8100 1595 8104 1648
rect 13427 1597 13436 1602
rect 8022 1590 8043 1594
rect 8034 1566 8040 1590
rect 8073 1566 8077 1588
rect 8144 1566 8149 1590
rect 12933 1571 12964 1574
rect 8034 1563 8153 1566
rect 12933 1526 12937 1571
rect 12960 1518 12964 1571
rect 12882 1513 12903 1517
rect 12894 1489 12900 1513
rect 12933 1489 12937 1511
rect 13004 1489 13009 1513
rect 12894 1486 13013 1489
rect 8078 1398 8109 1401
rect 8078 1353 8082 1398
rect 8105 1345 8109 1398
rect 12520 1398 12523 1404
rect 12520 1395 12557 1398
rect 12554 1392 12557 1395
rect 12554 1389 12575 1392
rect 12584 1376 12587 1386
rect 12521 1373 12587 1376
rect 8536 1353 8539 1359
rect 12521 1355 12524 1373
rect 8536 1350 8573 1353
rect 8570 1347 8573 1350
rect 8027 1340 8048 1344
rect 8039 1316 8045 1340
rect 8078 1316 8082 1338
rect 8149 1316 8154 1340
rect 8570 1344 8591 1347
rect 8600 1331 8603 1341
rect 8537 1328 8603 1331
rect 8039 1313 8158 1316
rect 8537 1310 8540 1328
rect 8076 1238 8107 1241
rect 8076 1193 8080 1238
rect 8103 1185 8107 1238
rect 8025 1180 8046 1184
rect 8037 1156 8043 1180
rect 8076 1156 8080 1178
rect 8147 1156 8152 1180
rect 8037 1153 8156 1156
rect 13478 1043 13487 1048
rect 12918 1018 12949 1021
rect 8529 1010 8532 1016
rect 8529 1007 8566 1010
rect 8104 1003 8135 1006
rect 8563 1004 8566 1007
rect 8104 958 8108 1003
rect 8131 950 8135 1003
rect 8563 1001 8584 1004
rect 8593 988 8596 998
rect 8530 985 8596 988
rect 8530 967 8533 985
rect 12460 968 12463 974
rect 12918 973 12922 1018
rect 12460 965 12497 968
rect 12945 965 12949 1018
rect 12494 962 12497 965
rect 12494 959 12515 962
rect 12867 960 12888 964
rect 8053 945 8074 949
rect 8065 921 8071 945
rect 12524 946 12527 956
rect 8104 921 8108 943
rect 8175 921 8180 945
rect 12461 943 12527 946
rect 12461 925 12464 943
rect 12879 936 12885 960
rect 12918 936 12922 958
rect 12989 936 12994 960
rect 12879 933 12998 936
rect 8065 918 8184 921
rect 8113 878 8144 881
rect 8113 833 8117 878
rect 8140 825 8144 878
rect 8062 820 8083 824
rect 8074 796 8080 820
rect 8113 796 8117 818
rect 8184 796 8189 820
rect 8074 793 8193 796
rect 12931 726 12962 729
rect 12931 681 12935 726
rect 12958 673 12962 726
rect 13463 694 13472 699
rect 12880 668 12901 672
rect 12892 644 12898 668
rect 12931 644 12935 666
rect 13002 644 13007 668
rect 12892 641 13011 644
rect 12417 432 12420 438
rect 12417 429 12454 432
rect 12451 426 12454 429
rect 12451 423 12472 426
rect 12481 410 12484 420
rect 12418 407 12484 410
rect 12418 389 12421 407
rect 12953 352 12984 355
rect 12953 307 12957 352
rect 12980 299 12984 352
rect 13516 309 13525 314
rect 12902 294 12923 298
rect 12914 270 12920 294
rect 12953 270 12957 292
rect 13024 270 13029 294
rect 12914 267 13033 270
<< m123contact >>
rect 12487 2245 12492 2250
rect 12487 2192 12492 2197
rect 12505 2196 12510 2201
rect 12519 2151 12524 2156
rect 8525 2108 8530 2113
rect 8525 2055 8530 2060
rect 8543 2059 8548 2064
rect 8557 2014 8562 2019
rect 8516 1749 8521 1754
rect 8516 1696 8521 1701
rect 8534 1700 8539 1705
rect 8548 1655 8553 1660
rect 12527 1435 12532 1440
rect 8543 1390 8548 1395
rect 12527 1382 12532 1387
rect 12545 1386 12550 1391
rect 8543 1337 8548 1342
rect 8561 1341 8566 1346
rect 12559 1341 12564 1346
rect 8575 1296 8580 1301
rect 8536 1047 8541 1052
rect 12467 1005 12472 1010
rect 8536 994 8541 999
rect 8554 998 8559 1003
rect 8568 953 8573 958
rect 12467 952 12472 957
rect 12485 956 12490 961
rect 12499 911 12504 916
rect 12424 469 12429 474
rect 12424 416 12429 421
rect 12442 420 12447 425
rect 12456 375 12461 380
<< metal3 >>
rect 12487 2197 12490 2245
rect 12510 2196 12522 2199
rect 12519 2156 12522 2196
rect 8525 2060 8528 2108
rect 8548 2059 8560 2062
rect 8557 2019 8560 2059
rect 8516 1701 8519 1749
rect 8539 1700 8551 1703
rect 8548 1660 8551 1700
rect 8543 1342 8546 1390
rect 12527 1387 12530 1435
rect 12550 1386 12562 1389
rect 12559 1346 12562 1386
rect 8566 1341 8578 1344
rect 8575 1301 8578 1341
rect 8536 999 8539 1047
rect 8559 998 8571 1001
rect 8568 958 8571 998
rect 12467 957 12470 1005
rect 12490 956 12502 959
rect 12499 916 12502 956
rect 12424 421 12427 469
rect 12447 420 12459 423
rect 12456 380 12459 420
<< labels >>
rlabel metal1 10165 1772 10169 1776 1 pdr1
rlabel metal2 10161 1656 10165 1661 2 prop_1
rlabel metal1 10173 1662 10177 1667 1 prop1_car0
rlabel metal1 10193 1771 10197 1776 1 prop1_car0
rlabel metal2 10189 1656 10193 1661 1 carry_0
rlabel metal1 10201 1662 10205 1667 1 clock_car0
rlabel metal1 10220 1771 10224 1776 1 clock_car0
rlabel metal2 10216 1656 10220 1661 1 clock_in
rlabel metal1 10228 1662 10232 1667 1 gnd!
rlabel metal1 10259 1771 10263 1776 1 pdr2
rlabel metal2 10255 1656 10259 1661 1 prop_2
rlabel metal1 10267 1662 10271 1667 1 pdr1
rlabel metal1 10287 1771 10291 1776 1 pdr1
rlabel metal2 10283 1656 10287 1661 1 gen_1
rlabel metal1 10295 1662 10299 1667 1 clock_car0
rlabel metal1 10314 1771 10318 1776 1 pdr3
rlabel metal2 10310 1656 10314 1661 1 prop_3
rlabel metal1 10322 1662 10326 1667 1 pdr2
rlabel metal1 10354 1772 10358 1777 1 pdr2
rlabel metal2 10350 1657 10354 1662 1 gen_2
rlabel metal1 10362 1663 10366 1668 1 clock_car0
rlabel metal1 10382 1772 10386 1777 1 pdr4
rlabel metal2 10378 1657 10382 1662 1 prop_4
rlabel metal1 10390 1663 10394 1668 1 pdr3
rlabel metal1 10409 1772 10413 1777 1 pdr3
rlabel metal2 10405 1657 10409 1662 1 gen_3
rlabel metal1 10417 1663 10421 1668 1 clock_car0
rlabel metal1 10445 1772 10449 1777 1 pdr4
rlabel metal2 10441 1657 10445 1662 1 gen_4
rlabel metal1 10453 1663 10457 1668 7 clock_car0
rlabel metal1 10229 2019 10233 2024 5 vdd!
rlabel metal1 10279 2020 10283 2025 5 vdd!
rlabel metal1 10329 2020 10333 2025 5 vdd!
rlabel metal1 10376 2020 10380 2025 5 vdd!
rlabel metal2 10218 1931 10224 1937 2 clock_in
rlabel metal2 10268 1932 10274 1938 1 clock_in
rlabel metal2 10318 1932 10324 1938 1 clock_in
rlabel metal2 10365 1932 10370 1938 1 clock_in
rlabel metal1 10237 1940 10241 1945 1 pdr1
rlabel metal1 10287 1941 10291 1945 1 pdr2
rlabel metal1 10337 1941 10341 1945 1 pdr3
rlabel metal1 10384 1941 10388 1945 1 pdr4
rlabel metal1 10823 1682 10827 1686 1 gnd!
rlabel metal1 10819 1786 10824 1790 5 vdd!
rlabel metal2 10695 1718 10698 1723 1 pdr1
rlabel metal2 10733 1718 10736 1723 1 pdr2
rlabel metal2 10777 1718 10780 1723 1 pdr3
rlabel metal2 10815 1718 10818 1723 1 pdr4
rlabel metal1 10706 1718 10710 1723 1 c1
rlabel metal1 10744 1718 10748 1723 1 c2
rlabel metal1 10788 1718 10792 1723 1 c3
rlabel metal1 10826 1718 10830 1723 1 c4
rlabel metal1 10869 1684 10873 1688 1 gnd!
rlabel metal1 10865 1788 10870 1792 5 vdd!
rlabel metal2 10861 1720 10864 1725 1 clk_org
rlabel metal1 10872 1720 10876 1725 1 clock_in
rlabel metal1 10698 1786 10702 1790 5 vdd!
rlabel metal1 10736 1786 10740 1790 5 vdd!
rlabel metal1 10780 1786 10784 1790 5 vdd!
rlabel metal1 10784 1682 10788 1686 1 gnd!
rlabel metal1 10747 1682 10751 1686 1 gnd!
rlabel metal1 10707 1682 10711 1686 1 gnd!
rlabel metal1 9028 1908 9028 1908 5 vdd
rlabel metal1 9029 1821 9029 1821 1 gnd
rlabel metal1 9061 1839 9061 1839 1 gnd
rlabel metal1 9058 1896 9058 1896 5 vdd
rlabel metal1 9030 1558 9030 1558 5 vdd
rlabel metal1 9031 1471 9031 1471 1 gnd
rlabel metal1 9063 1489 9063 1489 1 gnd
rlabel metal1 9060 1546 9060 1546 5 vdd
rlabel metal1 9038 1266 9038 1266 5 vdd
rlabel metal1 9039 1179 9039 1179 1 gnd
rlabel metal1 9071 1197 9071 1197 1 gnd
rlabel metal1 9068 1254 9068 1254 5 vdd
rlabel metal1 9026 900 9026 900 5 vdd
rlabel metal1 9027 813 9027 813 1 gnd
rlabel metal1 9059 831 9059 831 1 gnd
rlabel metal1 9056 888 9056 888 5 vdd
rlabel metal1 9013 1859 9013 1859 3 q_a1
rlabel metal1 9015 1852 9015 1852 3 q_b1
rlabel metal1 9077 1859 9077 1859 1 gen_1
rlabel metal1 9016 1508 9016 1508 1 q_a2
rlabel metal1 9016 1501 9016 1501 1 q_b2
rlabel metal1 9079 1510 9079 1510 1 gen_2
rlabel metal1 9023 1216 9023 1216 1 q_b3
rlabel metal1 9025 1209 9025 1209 1 q_a3
rlabel metal1 9086 1218 9086 1218 1 gen_3
rlabel metal1 9011 851 9011 851 3 q_a4
rlabel metal1 9011 845 9011 845 3 q_b4
rlabel metal1 9074 852 9074 852 1 gen_4
rlabel metal1 8543 2008 8547 2011 1 gnd
rlabel metal1 8593 2014 8596 2016 1 gnd
rlabel metal1 8541 2064 8542 2066 1 gnd
rlabel metal1 8537 2108 8540 2110 5 vdd
rlabel metal1 8538 2054 8541 2056 1 vdd
rlabel metal1 8534 1649 8538 1652 1 gnd
rlabel metal1 8584 1655 8587 1657 1 gnd
rlabel metal1 8532 1705 8533 1707 1 gnd
rlabel metal1 8528 1749 8531 1751 5 vdd
rlabel metal1 8529 1695 8532 1697 1 vdd
rlabel metal1 8561 1290 8565 1293 1 gnd
rlabel metal1 8611 1296 8614 1298 1 gnd
rlabel metal1 8559 1346 8560 1348 1 gnd
rlabel metal1 8555 1390 8558 1392 5 vdd
rlabel metal1 8556 1336 8559 1338 1 vdd
rlabel metal1 8554 947 8558 950 1 gnd
rlabel metal1 8604 953 8607 955 1 gnd
rlabel metal1 8552 1003 8553 1005 1 gnd
rlabel metal1 8548 1047 8551 1049 5 vdd
rlabel metal1 8549 993 8552 995 1 vdd
rlabel metal1 12505 2145 12509 2148 1 gnd
rlabel metal1 12555 2151 12558 2153 1 gnd
rlabel metal1 12503 2201 12504 2203 1 gnd
rlabel metal1 12499 2245 12502 2247 5 vdd
rlabel metal1 12500 2191 12503 2193 1 vdd
rlabel metal1 12545 1335 12549 1338 1 gnd
rlabel metal1 12595 1341 12598 1343 1 gnd
rlabel metal1 12543 1391 12544 1393 1 gnd
rlabel metal1 12539 1435 12542 1437 5 vdd
rlabel metal1 12540 1381 12543 1383 1 vdd
rlabel metal1 12485 905 12489 908 1 gnd
rlabel metal1 12535 911 12538 913 1 gnd
rlabel metal1 12483 961 12484 963 1 gnd
rlabel metal1 12479 1005 12482 1007 5 vdd
rlabel metal1 12480 951 12483 953 1 vdd
rlabel metal1 8515 2080 8515 2080 1 q_a1
rlabel metal1 8515 2026 8515 2026 1 q_b1
rlabel metal1 8631 2045 8631 2045 1 prop_1
rlabel metal1 8506 1721 8506 1721 3 q_a2
rlabel metal1 8506 1666 8506 1666 3 q_b2
rlabel metal1 8624 1687 8624 1687 1 prop_2
rlabel metal1 8534 1362 8534 1362 1 q_a3
rlabel metal1 8534 1308 8534 1308 1 q_b3
rlabel metal1 8651 1327 8651 1327 1 prop_3
rlabel metal1 8526 1018 8526 1018 1 q_a4
rlabel metal1 8526 965 8526 965 1 q_b4
rlabel metal1 8645 984 8645 984 1 prop_4
rlabel metal1 12477 2217 12477 2217 1 carry_0
rlabel metal1 12477 2163 12477 2163 1 prop_1
rlabel metal1 12596 2182 12596 2182 1 s1
rlabel metal1 12518 1406 12518 1406 1 c1
rlabel metal1 12517 1352 12517 1352 1 prop_2
rlabel metal1 12636 1371 12636 1371 7 s2
rlabel metal1 12457 977 12457 977 1 c2
rlabel metal1 12457 922 12457 922 1 prop_3
rlabel metal1 12576 942 12576 942 1 s3
rlabel metal1 12442 369 12446 372 1 gnd
rlabel metal1 12492 375 12495 377 1 gnd
rlabel metal1 12440 425 12441 427 1 gnd
rlabel metal1 12436 469 12439 471 5 vdd
rlabel metal1 12437 415 12440 417 1 vdd
rlabel metal1 12532 406 12532 406 1 s4
rlabel metal1 12414 387 12414 387 1 prop_4
rlabel metal1 12414 440 12414 440 1 c3
rlabel metal1 8000 2228 8003 2229 1 gnd
rlabel metal1 8006 2300 8008 2301 5 vdd
rlabel metal2 7987 2249 7987 2249 1 clk_org
rlabel metal1 8000 2048 8003 2049 1 gnd
rlabel metal1 8006 2120 8008 2121 5 vdd
rlabel metal2 7987 2069 7987 2069 1 clk_org
rlabel metal1 8006 2397 8009 2398 1 gnd
rlabel metal1 8012 2469 8014 2470 5 vdd
rlabel metal2 7993 2418 7993 2418 1 clk_org
rlabel metal1 8048 1732 8051 1733 1 gnd
rlabel metal1 8054 1804 8056 1805 5 vdd
rlabel metal2 8035 1753 8035 1753 1 clk_org
rlabel metal1 8052 1570 8055 1571 1 gnd
rlabel metal1 8058 1642 8060 1643 5 vdd
rlabel metal2 8039 1591 8039 1591 1 clk_org
rlabel metal1 8057 1320 8060 1321 1 gnd
rlabel metal1 8063 1392 8065 1393 5 vdd
rlabel metal2 8044 1341 8044 1341 1 clk_org
rlabel metal1 8055 1160 8058 1161 1 gnd
rlabel metal1 8061 1232 8063 1233 5 vdd
rlabel metal2 8042 1181 8042 1181 1 clk_org
rlabel metal1 8083 925 8086 926 1 gnd
rlabel metal1 8089 997 8091 998 5 vdd
rlabel metal2 8070 946 8070 946 1 clk_org
rlabel metal1 8092 800 8095 801 1 gnd
rlabel metal1 8098 872 8100 873 5 vdd
rlabel metal2 8079 821 8079 821 1 clk_org
rlabel metal1 7992 2427 7992 2427 1 cin
rlabel metal1 8149 2423 8149 2423 1 carry_0
rlabel metal1 7987 2258 7987 2258 1 a1
rlabel metal1 8142 2255 8142 2255 1 q_a1
rlabel metal1 7987 2078 7987 2078 1 b1
rlabel metal1 8142 2075 8142 2075 1 q_b1
rlabel metal1 8035 1762 8035 1762 1 a2
rlabel metal1 8190 1758 8190 1758 1 q_a2
rlabel metal1 8040 1600 8040 1600 1 b2
rlabel metal1 8193 1596 8193 1596 1 q_b2
rlabel metal1 8044 1350 8044 1350 1 a3
rlabel metal1 8198 1346 8198 1346 1 q_a3
rlabel metal1 8043 1190 8043 1190 1 b3
rlabel metal1 8198 1187 8198 1187 1 q_b3
rlabel metal1 8070 956 8070 956 1 a4
rlabel metal1 8225 951 8225 951 1 q_a4
rlabel metal1 8079 830 8079 830 1 b4
rlabel metal1 8234 827 8234 827 1 q_b4
rlabel metal1 12927 1934 12930 1935 1 gnd
rlabel metal1 12933 2006 12935 2007 5 vdd
rlabel metal2 12914 1955 12914 1955 1 clk_org
rlabel metal1 12912 1493 12915 1494 1 gnd
rlabel metal1 12918 1565 12920 1566 5 vdd
rlabel metal2 12899 1514 12899 1514 1 clk_org
rlabel metal1 12897 940 12900 941 1 gnd
rlabel metal1 12903 1012 12905 1013 5 vdd
rlabel metal2 12884 961 12884 961 1 clk_org
rlabel metal1 12910 648 12913 649 1 gnd
rlabel metal1 12916 720 12918 721 5 vdd
rlabel metal2 12897 669 12897 669 1 clk_org
rlabel metal1 12914 1964 12914 1964 1 s1
rlabel metal1 13069 1961 13069 1961 7 q_s1
rlabel metal1 12900 1523 12900 1523 1 s2
rlabel metal1 13053 1519 13053 1519 1 q_s2
rlabel metal1 12884 970 12884 970 1 s3
rlabel metal1 13039 967 13039 967 1 q_s3
rlabel metal1 12897 678 12897 678 1 s4
rlabel metal1 13051 674 13051 674 1 q_s4
rlabel metal1 12932 274 12935 275 1 gnd
rlabel metal1 12938 346 12940 347 5 vdd
rlabel metal2 12919 295 12919 295 1 clk_org
rlabel metal1 12919 304 12919 304 1 c4
rlabel metal1 13074 301 13074 301 7 q_c4
rlabel metal1 13411 2062 13411 2062 5 vdd!
rlabel metal1 13411 1998 13411 1998 1 gnd!
rlabel metal1 13439 1641 13439 1641 5 vdd!
rlabel metal1 13439 1577 13439 1577 1 gnd!
rlabel metal1 13490 1087 13490 1087 5 vdd!
rlabel metal1 13490 1023 13490 1023 1 gnd!
rlabel metal1 13475 738 13475 738 5 vdd!
rlabel metal1 13475 674 13475 674 1 gnd!
rlabel metal1 13528 353 13528 353 5 vdd!
rlabel metal1 13528 289 13528 289 1 gnd!
rlabel metal2 13401 2020 13401 2020 1 q_s1
rlabel metal1 13424 2021 13424 2021 1 iq_s1
rlabel metal2 13430 1599 13430 1599 1 q_s2
rlabel metal1 13451 1600 13451 1600 1 iq_s2
rlabel metal2 13480 1045 13480 1045 1 q_s3
rlabel metal1 13502 1046 13502 1046 1 iq_s3
rlabel metal2 13466 697 13466 697 1 q_s4
rlabel metal1 13487 697 13487 697 1 iq_s4
rlabel metal2 13518 312 13518 312 1 q_c4
rlabel metal1 13540 311 13540 311 7 iq_c4
<< end >>
