magic
tech scmos
timestamp 1732014888
<< nwell >>
rect -833 -1000 -801 -963
rect -795 -1000 -769 -963
rect -751 -1000 -725 -963
rect -706 -1000 -680 -963
rect -839 -1169 -807 -1132
rect -801 -1169 -775 -1132
rect -757 -1169 -731 -1132
rect -712 -1169 -686 -1132
rect 3658 -1209 3682 -1185
rect 3697 -1195 3731 -1189
rect 3697 -1225 3759 -1195
rect 3725 -1231 3759 -1225
rect 3658 -1264 3682 -1240
rect -839 -1349 -807 -1312
rect -801 -1349 -775 -1312
rect -757 -1349 -731 -1312
rect -712 -1349 -686 -1312
rect -304 -1346 -280 -1322
rect -265 -1332 -231 -1326
rect -265 -1362 -203 -1332
rect -237 -1368 -203 -1362
rect -304 -1401 -280 -1377
rect 1394 -1482 1418 -1420
rect 1444 -1481 1468 -1419
rect 1494 -1481 1518 -1419
rect 1541 -1481 1565 -1419
rect 4088 -1463 4120 -1426
rect 4126 -1463 4152 -1426
rect 4170 -1463 4196 -1426
rect 4215 -1463 4241 -1426
rect 183 -1560 219 -1520
rect 225 -1567 249 -1527
rect -791 -1665 -759 -1628
rect -753 -1665 -727 -1628
rect -709 -1665 -683 -1628
rect -664 -1665 -638 -1628
rect -313 -1705 -289 -1681
rect -274 -1691 -240 -1685
rect -274 -1721 -212 -1691
rect 1863 -1703 1887 -1651
rect 1901 -1703 1925 -1651
rect 1945 -1703 1969 -1651
rect 1983 -1703 2007 -1651
rect 2029 -1701 2053 -1649
rect -246 -1727 -212 -1721
rect -313 -1760 -289 -1736
rect -787 -1827 -755 -1790
rect -749 -1827 -723 -1790
rect -705 -1827 -679 -1790
rect -660 -1827 -634 -1790
rect 185 -1910 221 -1870
rect 227 -1917 251 -1877
rect 4073 -1904 4105 -1867
rect 4111 -1904 4137 -1867
rect 4155 -1904 4181 -1867
rect 4200 -1904 4226 -1867
rect 3698 -2019 3722 -1995
rect 3737 -2005 3771 -1999
rect 3737 -2035 3799 -2005
rect -782 -2077 -750 -2040
rect -744 -2077 -718 -2040
rect -700 -2077 -674 -2040
rect -655 -2077 -629 -2040
rect -286 -2064 -262 -2040
rect 3765 -2041 3799 -2035
rect -247 -2050 -213 -2044
rect -247 -2080 -185 -2050
rect 3698 -2074 3722 -2050
rect -219 -2086 -185 -2080
rect -286 -2119 -262 -2095
rect -784 -2237 -752 -2200
rect -746 -2237 -720 -2200
rect -702 -2237 -676 -2200
rect -657 -2237 -631 -2200
rect 193 -2202 229 -2162
rect 235 -2209 259 -2169
rect -293 -2407 -269 -2383
rect -254 -2393 -220 -2387
rect -254 -2423 -192 -2393
rect -226 -2429 -192 -2423
rect -756 -2472 -724 -2435
rect -718 -2472 -692 -2435
rect -674 -2472 -648 -2435
rect -629 -2472 -603 -2435
rect -293 -2462 -269 -2438
rect 3638 -2449 3662 -2425
rect 3677 -2435 3711 -2429
rect 3677 -2465 3739 -2435
rect 4058 -2457 4090 -2420
rect 4096 -2457 4122 -2420
rect 4140 -2457 4166 -2420
rect 4185 -2457 4211 -2420
rect 3705 -2471 3739 -2465
rect 3638 -2504 3662 -2480
rect -747 -2597 -715 -2560
rect -709 -2597 -683 -2560
rect -665 -2597 -639 -2560
rect -620 -2597 -594 -2560
rect 181 -2568 217 -2528
rect 223 -2575 247 -2535
rect 4071 -2749 4103 -2712
rect 4109 -2749 4135 -2712
rect 4153 -2749 4179 -2712
rect 4198 -2749 4224 -2712
rect 3595 -2985 3619 -2961
rect 3634 -2971 3668 -2965
rect 3634 -3001 3696 -2971
rect 3662 -3007 3696 -3001
rect 3595 -3040 3619 -3016
rect 4093 -3123 4125 -3086
rect 4131 -3123 4157 -3086
rect 4175 -3123 4201 -3086
rect 4220 -3123 4246 -3086
<< ntransistor >>
rect -826 -1026 -824 -1016
rect -790 -1026 -788 -1016
rect -782 -1026 -780 -1016
rect -746 -1026 -744 -1016
rect -738 -1026 -736 -1016
rect -695 -1026 -693 -1016
rect -832 -1195 -830 -1185
rect -796 -1195 -794 -1185
rect -788 -1195 -786 -1185
rect -752 -1195 -750 -1185
rect -744 -1195 -742 -1185
rect -701 -1195 -699 -1185
rect 3669 -1223 3671 -1217
rect 3708 -1272 3710 -1260
rect 3718 -1272 3720 -1260
rect 3736 -1272 3738 -1260
rect 3746 -1272 3748 -1260
rect 3669 -1278 3671 -1272
rect -293 -1360 -291 -1354
rect -832 -1375 -830 -1365
rect -796 -1375 -794 -1365
rect -788 -1375 -786 -1365
rect -752 -1375 -750 -1365
rect -744 -1375 -742 -1365
rect -701 -1375 -699 -1365
rect -254 -1409 -252 -1397
rect -244 -1409 -242 -1397
rect -226 -1409 -224 -1397
rect -216 -1409 -214 -1397
rect -293 -1415 -291 -1409
rect 4095 -1489 4097 -1479
rect 4131 -1489 4133 -1479
rect 4139 -1489 4141 -1479
rect 4175 -1489 4177 -1479
rect 4183 -1489 4185 -1479
rect 4226 -1489 4228 -1479
rect 194 -1603 196 -1583
rect 205 -1603 207 -1583
rect 236 -1585 238 -1575
rect -784 -1691 -782 -1681
rect -748 -1691 -746 -1681
rect -740 -1691 -738 -1681
rect -704 -1691 -702 -1681
rect -696 -1691 -694 -1681
rect -653 -1691 -651 -1681
rect -302 -1719 -300 -1713
rect -263 -1768 -261 -1756
rect -253 -1768 -251 -1756
rect -235 -1768 -233 -1756
rect -225 -1768 -223 -1756
rect 1341 -1762 1343 -1662
rect 1369 -1762 1371 -1662
rect 1396 -1762 1398 -1662
rect 1435 -1762 1437 -1662
rect 1463 -1762 1465 -1662
rect 1490 -1762 1492 -1662
rect 1530 -1761 1532 -1661
rect 1558 -1761 1560 -1661
rect 1585 -1761 1587 -1661
rect 1621 -1761 1623 -1661
rect 1874 -1735 1876 -1715
rect 1912 -1735 1914 -1715
rect 1956 -1735 1958 -1715
rect 1994 -1735 1996 -1715
rect 2040 -1733 2042 -1713
rect -302 -1774 -300 -1768
rect -780 -1853 -778 -1843
rect -744 -1853 -742 -1843
rect -736 -1853 -734 -1843
rect -700 -1853 -698 -1843
rect -692 -1853 -690 -1843
rect -649 -1853 -647 -1843
rect 196 -1953 198 -1933
rect 207 -1953 209 -1933
rect 238 -1935 240 -1925
rect 4080 -1930 4082 -1920
rect 4116 -1930 4118 -1920
rect 4124 -1930 4126 -1920
rect 4160 -1930 4162 -1920
rect 4168 -1930 4170 -1920
rect 4211 -1930 4213 -1920
rect 3709 -2033 3711 -2027
rect -275 -2078 -273 -2072
rect -775 -2103 -773 -2093
rect -739 -2103 -737 -2093
rect -731 -2103 -729 -2093
rect -695 -2103 -693 -2093
rect -687 -2103 -685 -2093
rect -644 -2103 -642 -2093
rect 3748 -2082 3750 -2070
rect 3758 -2082 3760 -2070
rect 3776 -2082 3778 -2070
rect 3786 -2082 3788 -2070
rect 3709 -2088 3711 -2082
rect -236 -2127 -234 -2115
rect -226 -2127 -224 -2115
rect -208 -2127 -206 -2115
rect -198 -2127 -196 -2115
rect -275 -2133 -273 -2127
rect 204 -2245 206 -2225
rect 215 -2245 217 -2225
rect 246 -2227 248 -2217
rect -777 -2263 -775 -2253
rect -741 -2263 -739 -2253
rect -733 -2263 -731 -2253
rect -697 -2263 -695 -2253
rect -689 -2263 -687 -2253
rect -646 -2263 -644 -2253
rect -282 -2421 -280 -2415
rect -243 -2470 -241 -2458
rect -233 -2470 -231 -2458
rect -215 -2470 -213 -2458
rect -205 -2470 -203 -2458
rect 3649 -2463 3651 -2457
rect -282 -2476 -280 -2470
rect -749 -2498 -747 -2488
rect -713 -2498 -711 -2488
rect -705 -2498 -703 -2488
rect -669 -2498 -667 -2488
rect -661 -2498 -659 -2488
rect -618 -2498 -616 -2488
rect 4065 -2483 4067 -2473
rect 4101 -2483 4103 -2473
rect 4109 -2483 4111 -2473
rect 4145 -2483 4147 -2473
rect 4153 -2483 4155 -2473
rect 4196 -2483 4198 -2473
rect 3688 -2512 3690 -2500
rect 3698 -2512 3700 -2500
rect 3716 -2512 3718 -2500
rect 3726 -2512 3728 -2500
rect 3649 -2518 3651 -2512
rect 192 -2611 194 -2591
rect 203 -2611 205 -2591
rect 234 -2593 236 -2583
rect -740 -2623 -738 -2613
rect -704 -2623 -702 -2613
rect -696 -2623 -694 -2613
rect -660 -2623 -658 -2613
rect -652 -2623 -650 -2613
rect -609 -2623 -607 -2613
rect 4078 -2775 4080 -2765
rect 4114 -2775 4116 -2765
rect 4122 -2775 4124 -2765
rect 4158 -2775 4160 -2765
rect 4166 -2775 4168 -2765
rect 4209 -2775 4211 -2765
rect 3606 -2999 3608 -2993
rect 3645 -3048 3647 -3036
rect 3655 -3048 3657 -3036
rect 3673 -3048 3675 -3036
rect 3683 -3048 3685 -3036
rect 3606 -3054 3608 -3048
rect 4100 -3149 4102 -3139
rect 4136 -3149 4138 -3139
rect 4144 -3149 4146 -3139
rect 4180 -3149 4182 -3139
rect 4188 -3149 4190 -3139
rect 4231 -3149 4233 -3139
<< ptransistor >>
rect -822 -994 -820 -969
rect -814 -994 -812 -969
rect -784 -994 -782 -969
rect -740 -994 -738 -969
rect -695 -994 -693 -969
rect -828 -1163 -826 -1138
rect -820 -1163 -818 -1138
rect -790 -1163 -788 -1138
rect -746 -1163 -744 -1138
rect -701 -1163 -699 -1138
rect 3669 -1203 3671 -1191
rect 3708 -1219 3710 -1195
rect 3718 -1219 3720 -1195
rect 3736 -1225 3738 -1201
rect 3746 -1225 3748 -1201
rect 3669 -1258 3671 -1246
rect -828 -1343 -826 -1318
rect -820 -1343 -818 -1318
rect -790 -1343 -788 -1318
rect -746 -1343 -744 -1318
rect -701 -1343 -699 -1318
rect -293 -1340 -291 -1328
rect -254 -1356 -252 -1332
rect -244 -1356 -242 -1332
rect -226 -1362 -224 -1338
rect -216 -1362 -214 -1338
rect -293 -1395 -291 -1383
rect 1405 -1476 1407 -1426
rect 1455 -1475 1457 -1425
rect 1505 -1475 1507 -1425
rect 1552 -1475 1554 -1425
rect 4099 -1457 4101 -1432
rect 4107 -1457 4109 -1432
rect 4137 -1457 4139 -1432
rect 4181 -1457 4183 -1432
rect 4226 -1457 4228 -1432
rect 194 -1554 196 -1534
rect 205 -1554 207 -1534
rect 236 -1561 238 -1541
rect -780 -1659 -778 -1634
rect -772 -1659 -770 -1634
rect -742 -1659 -740 -1634
rect -698 -1659 -696 -1634
rect -653 -1659 -651 -1634
rect -302 -1699 -300 -1687
rect -263 -1715 -261 -1691
rect -253 -1715 -251 -1691
rect -235 -1721 -233 -1697
rect -225 -1721 -223 -1697
rect -302 -1754 -300 -1742
rect 1874 -1697 1876 -1657
rect 1912 -1697 1914 -1657
rect 1956 -1697 1958 -1657
rect 1994 -1697 1996 -1657
rect 2040 -1695 2042 -1655
rect -776 -1821 -774 -1796
rect -768 -1821 -766 -1796
rect -738 -1821 -736 -1796
rect -694 -1821 -692 -1796
rect -649 -1821 -647 -1796
rect 196 -1904 198 -1884
rect 207 -1904 209 -1884
rect 238 -1911 240 -1891
rect 4084 -1898 4086 -1873
rect 4092 -1898 4094 -1873
rect 4122 -1898 4124 -1873
rect 4166 -1898 4168 -1873
rect 4211 -1898 4213 -1873
rect 3709 -2013 3711 -2001
rect 3748 -2029 3750 -2005
rect 3758 -2029 3760 -2005
rect 3776 -2035 3778 -2011
rect 3786 -2035 3788 -2011
rect -771 -2071 -769 -2046
rect -763 -2071 -761 -2046
rect -733 -2071 -731 -2046
rect -689 -2071 -687 -2046
rect -644 -2071 -642 -2046
rect -275 -2058 -273 -2046
rect -236 -2074 -234 -2050
rect -226 -2074 -224 -2050
rect -208 -2080 -206 -2056
rect -198 -2080 -196 -2056
rect 3709 -2068 3711 -2056
rect -275 -2113 -273 -2101
rect 204 -2196 206 -2176
rect 215 -2196 217 -2176
rect -773 -2231 -771 -2206
rect -765 -2231 -763 -2206
rect -735 -2231 -733 -2206
rect -691 -2231 -689 -2206
rect -646 -2231 -644 -2206
rect 246 -2203 248 -2183
rect -282 -2401 -280 -2389
rect -243 -2417 -241 -2393
rect -233 -2417 -231 -2393
rect -215 -2423 -213 -2399
rect -205 -2423 -203 -2399
rect -745 -2466 -743 -2441
rect -737 -2466 -735 -2441
rect -707 -2466 -705 -2441
rect -663 -2466 -661 -2441
rect -618 -2466 -616 -2441
rect -282 -2456 -280 -2444
rect 3649 -2443 3651 -2431
rect 3688 -2459 3690 -2435
rect 3698 -2459 3700 -2435
rect 3716 -2465 3718 -2441
rect 3726 -2465 3728 -2441
rect 4069 -2451 4071 -2426
rect 4077 -2451 4079 -2426
rect 4107 -2451 4109 -2426
rect 4151 -2451 4153 -2426
rect 4196 -2451 4198 -2426
rect 3649 -2498 3651 -2486
rect 192 -2562 194 -2542
rect 203 -2562 205 -2542
rect -736 -2591 -734 -2566
rect -728 -2591 -726 -2566
rect -698 -2591 -696 -2566
rect -654 -2591 -652 -2566
rect -609 -2591 -607 -2566
rect 234 -2569 236 -2549
rect 4082 -2743 4084 -2718
rect 4090 -2743 4092 -2718
rect 4120 -2743 4122 -2718
rect 4164 -2743 4166 -2718
rect 4209 -2743 4211 -2718
rect 3606 -2979 3608 -2967
rect 3645 -2995 3647 -2971
rect 3655 -2995 3657 -2971
rect 3673 -3001 3675 -2977
rect 3683 -3001 3685 -2977
rect 3606 -3034 3608 -3022
rect 4104 -3117 4106 -3092
rect 4112 -3117 4114 -3092
rect 4142 -3117 4144 -3092
rect 4186 -3117 4188 -3092
rect 4231 -3117 4233 -3092
<< ndiffusion >>
rect -827 -1026 -826 -1016
rect -824 -1026 -823 -1016
rect -791 -1026 -790 -1016
rect -788 -1026 -787 -1016
rect -783 -1026 -782 -1016
rect -780 -1026 -779 -1016
rect -747 -1026 -746 -1016
rect -744 -1026 -743 -1016
rect -739 -1026 -738 -1016
rect -736 -1026 -735 -1016
rect -696 -1026 -695 -1016
rect -693 -1026 -692 -1016
rect -833 -1195 -832 -1185
rect -830 -1195 -829 -1185
rect -797 -1195 -796 -1185
rect -794 -1195 -793 -1185
rect -789 -1195 -788 -1185
rect -786 -1195 -785 -1185
rect -753 -1195 -752 -1185
rect -750 -1195 -749 -1185
rect -745 -1195 -744 -1185
rect -742 -1195 -741 -1185
rect -702 -1195 -701 -1185
rect -699 -1195 -698 -1185
rect 3668 -1223 3669 -1217
rect 3671 -1223 3672 -1217
rect 3707 -1272 3708 -1260
rect 3710 -1272 3718 -1260
rect 3720 -1272 3721 -1260
rect 3735 -1272 3736 -1260
rect 3738 -1272 3746 -1260
rect 3748 -1272 3749 -1260
rect 3668 -1278 3669 -1272
rect 3671 -1278 3672 -1272
rect -294 -1360 -293 -1354
rect -291 -1360 -290 -1354
rect -833 -1375 -832 -1365
rect -830 -1375 -829 -1365
rect -797 -1375 -796 -1365
rect -794 -1375 -793 -1365
rect -789 -1375 -788 -1365
rect -786 -1375 -785 -1365
rect -753 -1375 -752 -1365
rect -750 -1375 -749 -1365
rect -745 -1375 -744 -1365
rect -742 -1375 -741 -1365
rect -702 -1375 -701 -1365
rect -699 -1375 -698 -1365
rect -255 -1409 -254 -1397
rect -252 -1409 -244 -1397
rect -242 -1409 -241 -1397
rect -227 -1409 -226 -1397
rect -224 -1409 -216 -1397
rect -214 -1409 -213 -1397
rect -294 -1415 -293 -1409
rect -291 -1415 -290 -1409
rect 4094 -1489 4095 -1479
rect 4097 -1489 4098 -1479
rect 4130 -1489 4131 -1479
rect 4133 -1489 4134 -1479
rect 4138 -1489 4139 -1479
rect 4141 -1489 4142 -1479
rect 4174 -1489 4175 -1479
rect 4177 -1489 4178 -1479
rect 4182 -1489 4183 -1479
rect 4185 -1489 4186 -1479
rect 4225 -1489 4226 -1479
rect 4228 -1489 4229 -1479
rect 193 -1603 194 -1583
rect 196 -1603 205 -1583
rect 207 -1603 208 -1583
rect 235 -1585 236 -1575
rect 238 -1585 239 -1575
rect -785 -1691 -784 -1681
rect -782 -1691 -781 -1681
rect -749 -1691 -748 -1681
rect -746 -1691 -745 -1681
rect -741 -1691 -740 -1681
rect -738 -1691 -737 -1681
rect -705 -1691 -704 -1681
rect -702 -1691 -701 -1681
rect -697 -1691 -696 -1681
rect -694 -1691 -693 -1681
rect -654 -1691 -653 -1681
rect -651 -1691 -650 -1681
rect -303 -1719 -302 -1713
rect -300 -1719 -299 -1713
rect -264 -1768 -263 -1756
rect -261 -1768 -253 -1756
rect -251 -1768 -250 -1756
rect -236 -1768 -235 -1756
rect -233 -1768 -225 -1756
rect -223 -1768 -222 -1756
rect 1340 -1762 1341 -1662
rect 1343 -1762 1344 -1662
rect 1368 -1762 1369 -1662
rect 1371 -1762 1372 -1662
rect 1395 -1762 1396 -1662
rect 1398 -1762 1399 -1662
rect 1434 -1762 1435 -1662
rect 1437 -1762 1438 -1662
rect 1462 -1762 1463 -1662
rect 1465 -1762 1466 -1662
rect 1489 -1762 1490 -1662
rect 1492 -1762 1493 -1662
rect 1529 -1761 1530 -1661
rect 1532 -1761 1533 -1661
rect 1557 -1761 1558 -1661
rect 1560 -1761 1561 -1661
rect 1584 -1761 1585 -1661
rect 1587 -1761 1588 -1661
rect 1620 -1761 1621 -1661
rect 1623 -1761 1624 -1661
rect 1873 -1735 1874 -1715
rect 1876 -1735 1877 -1715
rect 1911 -1735 1912 -1715
rect 1914 -1735 1915 -1715
rect 1955 -1735 1956 -1715
rect 1958 -1735 1959 -1715
rect 1993 -1735 1994 -1715
rect 1996 -1735 1997 -1715
rect 2039 -1733 2040 -1713
rect 2042 -1733 2043 -1713
rect -303 -1774 -302 -1768
rect -300 -1774 -299 -1768
rect -781 -1853 -780 -1843
rect -778 -1853 -777 -1843
rect -745 -1853 -744 -1843
rect -742 -1853 -741 -1843
rect -737 -1853 -736 -1843
rect -734 -1853 -733 -1843
rect -701 -1853 -700 -1843
rect -698 -1853 -697 -1843
rect -693 -1853 -692 -1843
rect -690 -1853 -689 -1843
rect -650 -1853 -649 -1843
rect -647 -1853 -646 -1843
rect 195 -1953 196 -1933
rect 198 -1953 207 -1933
rect 209 -1953 210 -1933
rect 237 -1935 238 -1925
rect 240 -1935 241 -1925
rect 4079 -1930 4080 -1920
rect 4082 -1930 4083 -1920
rect 4115 -1930 4116 -1920
rect 4118 -1930 4119 -1920
rect 4123 -1930 4124 -1920
rect 4126 -1930 4127 -1920
rect 4159 -1930 4160 -1920
rect 4162 -1930 4163 -1920
rect 4167 -1930 4168 -1920
rect 4170 -1930 4171 -1920
rect 4210 -1930 4211 -1920
rect 4213 -1930 4214 -1920
rect 3708 -2033 3709 -2027
rect 3711 -2033 3712 -2027
rect -276 -2078 -275 -2072
rect -273 -2078 -272 -2072
rect -776 -2103 -775 -2093
rect -773 -2103 -772 -2093
rect -740 -2103 -739 -2093
rect -737 -2103 -736 -2093
rect -732 -2103 -731 -2093
rect -729 -2103 -728 -2093
rect -696 -2103 -695 -2093
rect -693 -2103 -692 -2093
rect -688 -2103 -687 -2093
rect -685 -2103 -684 -2093
rect -645 -2103 -644 -2093
rect -642 -2103 -641 -2093
rect 3747 -2082 3748 -2070
rect 3750 -2082 3758 -2070
rect 3760 -2082 3761 -2070
rect 3775 -2082 3776 -2070
rect 3778 -2082 3786 -2070
rect 3788 -2082 3789 -2070
rect 3708 -2088 3709 -2082
rect 3711 -2088 3712 -2082
rect -237 -2127 -236 -2115
rect -234 -2127 -226 -2115
rect -224 -2127 -223 -2115
rect -209 -2127 -208 -2115
rect -206 -2127 -198 -2115
rect -196 -2127 -195 -2115
rect -276 -2133 -275 -2127
rect -273 -2133 -272 -2127
rect 203 -2245 204 -2225
rect 206 -2245 215 -2225
rect 217 -2245 218 -2225
rect 245 -2227 246 -2217
rect 248 -2227 249 -2217
rect -778 -2263 -777 -2253
rect -775 -2263 -774 -2253
rect -742 -2263 -741 -2253
rect -739 -2263 -738 -2253
rect -734 -2263 -733 -2253
rect -731 -2263 -730 -2253
rect -698 -2263 -697 -2253
rect -695 -2263 -694 -2253
rect -690 -2263 -689 -2253
rect -687 -2263 -686 -2253
rect -647 -2263 -646 -2253
rect -644 -2263 -643 -2253
rect -283 -2421 -282 -2415
rect -280 -2421 -279 -2415
rect -244 -2470 -243 -2458
rect -241 -2470 -233 -2458
rect -231 -2470 -230 -2458
rect -216 -2470 -215 -2458
rect -213 -2470 -205 -2458
rect -203 -2470 -202 -2458
rect 3648 -2463 3649 -2457
rect 3651 -2463 3652 -2457
rect -283 -2476 -282 -2470
rect -280 -2476 -279 -2470
rect -750 -2498 -749 -2488
rect -747 -2498 -746 -2488
rect -714 -2498 -713 -2488
rect -711 -2498 -710 -2488
rect -706 -2498 -705 -2488
rect -703 -2498 -702 -2488
rect -670 -2498 -669 -2488
rect -667 -2498 -666 -2488
rect -662 -2498 -661 -2488
rect -659 -2498 -658 -2488
rect -619 -2498 -618 -2488
rect -616 -2498 -615 -2488
rect 4064 -2483 4065 -2473
rect 4067 -2483 4068 -2473
rect 4100 -2483 4101 -2473
rect 4103 -2483 4104 -2473
rect 4108 -2483 4109 -2473
rect 4111 -2483 4112 -2473
rect 4144 -2483 4145 -2473
rect 4147 -2483 4148 -2473
rect 4152 -2483 4153 -2473
rect 4155 -2483 4156 -2473
rect 4195 -2483 4196 -2473
rect 4198 -2483 4199 -2473
rect 3687 -2512 3688 -2500
rect 3690 -2512 3698 -2500
rect 3700 -2512 3701 -2500
rect 3715 -2512 3716 -2500
rect 3718 -2512 3726 -2500
rect 3728 -2512 3729 -2500
rect 3648 -2518 3649 -2512
rect 3651 -2518 3652 -2512
rect 191 -2611 192 -2591
rect 194 -2611 203 -2591
rect 205 -2611 206 -2591
rect 233 -2593 234 -2583
rect 236 -2593 237 -2583
rect -741 -2623 -740 -2613
rect -738 -2623 -737 -2613
rect -705 -2623 -704 -2613
rect -702 -2623 -701 -2613
rect -697 -2623 -696 -2613
rect -694 -2623 -693 -2613
rect -661 -2623 -660 -2613
rect -658 -2623 -657 -2613
rect -653 -2623 -652 -2613
rect -650 -2623 -649 -2613
rect -610 -2623 -609 -2613
rect -607 -2623 -606 -2613
rect 4077 -2775 4078 -2765
rect 4080 -2775 4081 -2765
rect 4113 -2775 4114 -2765
rect 4116 -2775 4117 -2765
rect 4121 -2775 4122 -2765
rect 4124 -2775 4125 -2765
rect 4157 -2775 4158 -2765
rect 4160 -2775 4161 -2765
rect 4165 -2775 4166 -2765
rect 4168 -2775 4169 -2765
rect 4208 -2775 4209 -2765
rect 4211 -2775 4212 -2765
rect 3605 -2999 3606 -2993
rect 3608 -2999 3609 -2993
rect 3644 -3048 3645 -3036
rect 3647 -3048 3655 -3036
rect 3657 -3048 3658 -3036
rect 3672 -3048 3673 -3036
rect 3675 -3048 3683 -3036
rect 3685 -3048 3686 -3036
rect 3605 -3054 3606 -3048
rect 3608 -3054 3609 -3048
rect 4099 -3149 4100 -3139
rect 4102 -3149 4103 -3139
rect 4135 -3149 4136 -3139
rect 4138 -3149 4139 -3139
rect 4143 -3149 4144 -3139
rect 4146 -3149 4147 -3139
rect 4179 -3149 4180 -3139
rect 4182 -3149 4183 -3139
rect 4187 -3149 4188 -3139
rect 4190 -3149 4191 -3139
rect 4230 -3149 4231 -3139
rect 4233 -3149 4234 -3139
<< pdiffusion >>
rect -823 -994 -822 -969
rect -820 -994 -819 -969
rect -815 -994 -814 -969
rect -812 -994 -811 -969
rect -785 -994 -784 -969
rect -782 -994 -781 -969
rect -741 -994 -740 -969
rect -738 -994 -737 -969
rect -696 -994 -695 -969
rect -693 -994 -692 -969
rect -829 -1163 -828 -1138
rect -826 -1163 -825 -1138
rect -821 -1163 -820 -1138
rect -818 -1163 -817 -1138
rect -791 -1163 -790 -1138
rect -788 -1163 -787 -1138
rect -747 -1163 -746 -1138
rect -744 -1163 -743 -1138
rect -702 -1163 -701 -1138
rect -699 -1163 -698 -1138
rect 3668 -1203 3669 -1191
rect 3671 -1203 3672 -1191
rect 3707 -1219 3708 -1195
rect 3710 -1219 3712 -1195
rect 3716 -1219 3718 -1195
rect 3720 -1219 3721 -1195
rect 3735 -1225 3736 -1201
rect 3738 -1225 3740 -1201
rect 3744 -1225 3746 -1201
rect 3748 -1225 3749 -1201
rect 3668 -1258 3669 -1246
rect 3671 -1258 3672 -1246
rect -829 -1343 -828 -1318
rect -826 -1343 -825 -1318
rect -821 -1343 -820 -1318
rect -818 -1343 -817 -1318
rect -791 -1343 -790 -1318
rect -788 -1343 -787 -1318
rect -747 -1343 -746 -1318
rect -744 -1343 -743 -1318
rect -702 -1343 -701 -1318
rect -699 -1343 -698 -1318
rect -294 -1340 -293 -1328
rect -291 -1340 -290 -1328
rect -255 -1356 -254 -1332
rect -252 -1356 -250 -1332
rect -246 -1356 -244 -1332
rect -242 -1356 -241 -1332
rect -227 -1362 -226 -1338
rect -224 -1362 -222 -1338
rect -218 -1362 -216 -1338
rect -214 -1362 -213 -1338
rect -294 -1395 -293 -1383
rect -291 -1395 -290 -1383
rect 1404 -1476 1405 -1426
rect 1407 -1476 1408 -1426
rect 1454 -1475 1455 -1425
rect 1457 -1475 1458 -1425
rect 1504 -1475 1505 -1425
rect 1507 -1475 1508 -1425
rect 1551 -1475 1552 -1425
rect 1554 -1475 1555 -1425
rect 4098 -1457 4099 -1432
rect 4101 -1457 4102 -1432
rect 4106 -1457 4107 -1432
rect 4109 -1457 4110 -1432
rect 4136 -1457 4137 -1432
rect 4139 -1457 4140 -1432
rect 4180 -1457 4181 -1432
rect 4183 -1457 4184 -1432
rect 4225 -1457 4226 -1432
rect 4228 -1457 4229 -1432
rect 193 -1554 194 -1534
rect 196 -1554 200 -1534
rect 204 -1554 205 -1534
rect 207 -1554 208 -1534
rect 235 -1561 236 -1541
rect 238 -1561 239 -1541
rect -781 -1659 -780 -1634
rect -778 -1659 -777 -1634
rect -773 -1659 -772 -1634
rect -770 -1659 -769 -1634
rect -743 -1659 -742 -1634
rect -740 -1659 -739 -1634
rect -699 -1659 -698 -1634
rect -696 -1659 -695 -1634
rect -654 -1659 -653 -1634
rect -651 -1659 -650 -1634
rect -303 -1699 -302 -1687
rect -300 -1699 -299 -1687
rect -264 -1715 -263 -1691
rect -261 -1715 -259 -1691
rect -255 -1715 -253 -1691
rect -251 -1715 -250 -1691
rect -236 -1721 -235 -1697
rect -233 -1721 -231 -1697
rect -227 -1721 -225 -1697
rect -223 -1721 -222 -1697
rect -303 -1754 -302 -1742
rect -300 -1754 -299 -1742
rect 1873 -1697 1874 -1657
rect 1876 -1697 1877 -1657
rect 1911 -1697 1912 -1657
rect 1914 -1697 1915 -1657
rect 1955 -1697 1956 -1657
rect 1958 -1697 1959 -1657
rect 1993 -1697 1994 -1657
rect 1996 -1697 1997 -1657
rect 2039 -1695 2040 -1655
rect 2042 -1695 2043 -1655
rect -777 -1821 -776 -1796
rect -774 -1821 -773 -1796
rect -769 -1821 -768 -1796
rect -766 -1821 -765 -1796
rect -739 -1821 -738 -1796
rect -736 -1821 -735 -1796
rect -695 -1821 -694 -1796
rect -692 -1821 -691 -1796
rect -650 -1821 -649 -1796
rect -647 -1821 -646 -1796
rect 195 -1904 196 -1884
rect 198 -1904 202 -1884
rect 206 -1904 207 -1884
rect 209 -1904 210 -1884
rect 237 -1911 238 -1891
rect 240 -1911 241 -1891
rect 4083 -1898 4084 -1873
rect 4086 -1898 4087 -1873
rect 4091 -1898 4092 -1873
rect 4094 -1898 4095 -1873
rect 4121 -1898 4122 -1873
rect 4124 -1898 4125 -1873
rect 4165 -1898 4166 -1873
rect 4168 -1898 4169 -1873
rect 4210 -1898 4211 -1873
rect 4213 -1898 4214 -1873
rect 3708 -2013 3709 -2001
rect 3711 -2013 3712 -2001
rect 3747 -2029 3748 -2005
rect 3750 -2029 3752 -2005
rect 3756 -2029 3758 -2005
rect 3760 -2029 3761 -2005
rect 3775 -2035 3776 -2011
rect 3778 -2035 3780 -2011
rect 3784 -2035 3786 -2011
rect 3788 -2035 3789 -2011
rect -772 -2071 -771 -2046
rect -769 -2071 -768 -2046
rect -764 -2071 -763 -2046
rect -761 -2071 -760 -2046
rect -734 -2071 -733 -2046
rect -731 -2071 -730 -2046
rect -690 -2071 -689 -2046
rect -687 -2071 -686 -2046
rect -645 -2071 -644 -2046
rect -642 -2071 -641 -2046
rect -276 -2058 -275 -2046
rect -273 -2058 -272 -2046
rect -237 -2074 -236 -2050
rect -234 -2074 -232 -2050
rect -228 -2074 -226 -2050
rect -224 -2074 -223 -2050
rect -209 -2080 -208 -2056
rect -206 -2080 -204 -2056
rect -200 -2080 -198 -2056
rect -196 -2080 -195 -2056
rect 3708 -2068 3709 -2056
rect 3711 -2068 3712 -2056
rect -276 -2113 -275 -2101
rect -273 -2113 -272 -2101
rect 203 -2196 204 -2176
rect 206 -2196 210 -2176
rect 214 -2196 215 -2176
rect 217 -2196 218 -2176
rect -774 -2231 -773 -2206
rect -771 -2231 -770 -2206
rect -766 -2231 -765 -2206
rect -763 -2231 -762 -2206
rect -736 -2231 -735 -2206
rect -733 -2231 -732 -2206
rect -692 -2231 -691 -2206
rect -689 -2231 -688 -2206
rect -647 -2231 -646 -2206
rect -644 -2231 -643 -2206
rect 245 -2203 246 -2183
rect 248 -2203 249 -2183
rect -283 -2401 -282 -2389
rect -280 -2401 -279 -2389
rect -244 -2417 -243 -2393
rect -241 -2417 -239 -2393
rect -235 -2417 -233 -2393
rect -231 -2417 -230 -2393
rect -216 -2423 -215 -2399
rect -213 -2423 -211 -2399
rect -207 -2423 -205 -2399
rect -203 -2423 -202 -2399
rect -746 -2466 -745 -2441
rect -743 -2466 -742 -2441
rect -738 -2466 -737 -2441
rect -735 -2466 -734 -2441
rect -708 -2466 -707 -2441
rect -705 -2466 -704 -2441
rect -664 -2466 -663 -2441
rect -661 -2466 -660 -2441
rect -619 -2466 -618 -2441
rect -616 -2466 -615 -2441
rect -283 -2456 -282 -2444
rect -280 -2456 -279 -2444
rect 3648 -2443 3649 -2431
rect 3651 -2443 3652 -2431
rect 3687 -2459 3688 -2435
rect 3690 -2459 3692 -2435
rect 3696 -2459 3698 -2435
rect 3700 -2459 3701 -2435
rect 3715 -2465 3716 -2441
rect 3718 -2465 3720 -2441
rect 3724 -2465 3726 -2441
rect 3728 -2465 3729 -2441
rect 4068 -2451 4069 -2426
rect 4071 -2451 4072 -2426
rect 4076 -2451 4077 -2426
rect 4079 -2451 4080 -2426
rect 4106 -2451 4107 -2426
rect 4109 -2451 4110 -2426
rect 4150 -2451 4151 -2426
rect 4153 -2451 4154 -2426
rect 4195 -2451 4196 -2426
rect 4198 -2451 4199 -2426
rect 3648 -2498 3649 -2486
rect 3651 -2498 3652 -2486
rect 191 -2562 192 -2542
rect 194 -2562 198 -2542
rect 202 -2562 203 -2542
rect 205 -2562 206 -2542
rect -737 -2591 -736 -2566
rect -734 -2591 -733 -2566
rect -729 -2591 -728 -2566
rect -726 -2591 -725 -2566
rect -699 -2591 -698 -2566
rect -696 -2591 -695 -2566
rect -655 -2591 -654 -2566
rect -652 -2591 -651 -2566
rect -610 -2591 -609 -2566
rect -607 -2591 -606 -2566
rect 233 -2569 234 -2549
rect 236 -2569 237 -2549
rect 4081 -2743 4082 -2718
rect 4084 -2743 4085 -2718
rect 4089 -2743 4090 -2718
rect 4092 -2743 4093 -2718
rect 4119 -2743 4120 -2718
rect 4122 -2743 4123 -2718
rect 4163 -2743 4164 -2718
rect 4166 -2743 4167 -2718
rect 4208 -2743 4209 -2718
rect 4211 -2743 4212 -2718
rect 3605 -2979 3606 -2967
rect 3608 -2979 3609 -2967
rect 3644 -2995 3645 -2971
rect 3647 -2995 3649 -2971
rect 3653 -2995 3655 -2971
rect 3657 -2995 3658 -2971
rect 3672 -3001 3673 -2977
rect 3675 -3001 3677 -2977
rect 3681 -3001 3683 -2977
rect 3685 -3001 3686 -2977
rect 3605 -3034 3606 -3022
rect 3608 -3034 3609 -3022
rect 4103 -3117 4104 -3092
rect 4106 -3117 4107 -3092
rect 4111 -3117 4112 -3092
rect 4114 -3117 4115 -3092
rect 4141 -3117 4142 -3092
rect 4144 -3117 4145 -3092
rect 4185 -3117 4186 -3092
rect 4188 -3117 4189 -3092
rect 4230 -3117 4231 -3092
rect 4233 -3117 4234 -3092
<< ndcontact >>
rect -831 -1026 -827 -1016
rect -823 -1026 -819 -1016
rect -795 -1026 -791 -1016
rect -787 -1026 -783 -1016
rect -779 -1026 -775 -1016
rect -751 -1026 -747 -1016
rect -743 -1026 -739 -1016
rect -735 -1026 -731 -1016
rect -700 -1026 -696 -1016
rect -692 -1026 -688 -1016
rect -837 -1195 -833 -1185
rect -829 -1195 -825 -1185
rect -801 -1195 -797 -1185
rect -793 -1195 -789 -1185
rect -785 -1195 -781 -1185
rect -757 -1195 -753 -1185
rect -749 -1195 -745 -1185
rect -741 -1195 -737 -1185
rect -706 -1195 -702 -1185
rect -698 -1195 -694 -1185
rect 3664 -1223 3668 -1217
rect 3672 -1223 3676 -1217
rect 3703 -1272 3707 -1260
rect 3721 -1272 3725 -1260
rect 3731 -1272 3735 -1260
rect 3749 -1272 3753 -1260
rect 3664 -1278 3668 -1272
rect 3672 -1278 3676 -1272
rect -298 -1360 -294 -1354
rect -290 -1360 -286 -1354
rect -837 -1375 -833 -1365
rect -829 -1375 -825 -1365
rect -801 -1375 -797 -1365
rect -793 -1375 -789 -1365
rect -785 -1375 -781 -1365
rect -757 -1375 -753 -1365
rect -749 -1375 -745 -1365
rect -741 -1375 -737 -1365
rect -706 -1375 -702 -1365
rect -698 -1375 -694 -1365
rect -259 -1409 -255 -1397
rect -241 -1409 -237 -1397
rect -231 -1409 -227 -1397
rect -213 -1409 -209 -1397
rect -298 -1415 -294 -1409
rect -290 -1415 -286 -1409
rect 4090 -1489 4094 -1479
rect 4098 -1489 4102 -1479
rect 4126 -1489 4130 -1479
rect 4134 -1489 4138 -1479
rect 4142 -1489 4146 -1479
rect 4170 -1489 4174 -1479
rect 4178 -1489 4182 -1479
rect 4186 -1489 4190 -1479
rect 4221 -1489 4225 -1479
rect 4229 -1489 4233 -1479
rect 189 -1603 193 -1583
rect 208 -1603 212 -1583
rect 231 -1585 235 -1575
rect 239 -1585 243 -1575
rect -789 -1691 -785 -1681
rect -781 -1691 -777 -1681
rect -753 -1691 -749 -1681
rect -745 -1691 -741 -1681
rect -737 -1691 -733 -1681
rect -709 -1691 -705 -1681
rect -701 -1691 -697 -1681
rect -693 -1691 -689 -1681
rect -658 -1691 -654 -1681
rect -650 -1691 -646 -1681
rect -307 -1719 -303 -1713
rect -299 -1719 -295 -1713
rect -268 -1768 -264 -1756
rect -250 -1768 -246 -1756
rect -240 -1768 -236 -1756
rect -222 -1768 -218 -1756
rect 1336 -1762 1340 -1662
rect 1344 -1762 1348 -1662
rect 1364 -1762 1368 -1662
rect 1372 -1762 1376 -1662
rect 1391 -1762 1395 -1662
rect 1399 -1762 1403 -1662
rect 1430 -1762 1434 -1662
rect 1438 -1762 1442 -1662
rect 1458 -1762 1462 -1662
rect 1466 -1762 1470 -1662
rect 1485 -1762 1489 -1662
rect 1493 -1762 1497 -1662
rect 1525 -1761 1529 -1661
rect 1533 -1761 1537 -1661
rect 1553 -1761 1557 -1661
rect 1561 -1761 1565 -1661
rect 1580 -1761 1584 -1661
rect 1588 -1761 1592 -1661
rect 1616 -1761 1620 -1661
rect 1624 -1761 1628 -1661
rect 1869 -1735 1873 -1715
rect 1877 -1735 1881 -1715
rect 1907 -1735 1911 -1715
rect 1915 -1735 1919 -1715
rect 1951 -1735 1955 -1715
rect 1959 -1735 1963 -1715
rect 1989 -1735 1993 -1715
rect 1997 -1735 2001 -1715
rect 2035 -1733 2039 -1713
rect 2043 -1733 2047 -1713
rect -307 -1774 -303 -1768
rect -299 -1774 -295 -1768
rect -785 -1853 -781 -1843
rect -777 -1853 -773 -1843
rect -749 -1853 -745 -1843
rect -741 -1853 -737 -1843
rect -733 -1853 -729 -1843
rect -705 -1853 -701 -1843
rect -697 -1853 -693 -1843
rect -689 -1853 -685 -1843
rect -654 -1853 -650 -1843
rect -646 -1853 -642 -1843
rect 191 -1953 195 -1933
rect 210 -1953 214 -1933
rect 233 -1935 237 -1925
rect 241 -1935 245 -1925
rect 4075 -1930 4079 -1920
rect 4083 -1930 4087 -1920
rect 4111 -1930 4115 -1920
rect 4119 -1930 4123 -1920
rect 4127 -1930 4131 -1920
rect 4155 -1930 4159 -1920
rect 4163 -1930 4167 -1920
rect 4171 -1930 4175 -1920
rect 4206 -1930 4210 -1920
rect 4214 -1930 4218 -1920
rect 3704 -2033 3708 -2027
rect 3712 -2033 3716 -2027
rect -280 -2078 -276 -2072
rect -272 -2078 -268 -2072
rect -780 -2103 -776 -2093
rect -772 -2103 -768 -2093
rect -744 -2103 -740 -2093
rect -736 -2103 -732 -2093
rect -728 -2103 -724 -2093
rect -700 -2103 -696 -2093
rect -692 -2103 -688 -2093
rect -684 -2103 -680 -2093
rect -649 -2103 -645 -2093
rect -641 -2103 -637 -2093
rect 3743 -2082 3747 -2070
rect 3761 -2082 3765 -2070
rect 3771 -2082 3775 -2070
rect 3789 -2082 3793 -2070
rect 3704 -2088 3708 -2082
rect 3712 -2088 3716 -2082
rect -241 -2127 -237 -2115
rect -223 -2127 -219 -2115
rect -213 -2127 -209 -2115
rect -195 -2127 -191 -2115
rect -280 -2133 -276 -2127
rect -272 -2133 -268 -2127
rect 199 -2245 203 -2225
rect 218 -2245 222 -2225
rect 241 -2227 245 -2217
rect 249 -2227 253 -2217
rect -782 -2263 -778 -2253
rect -774 -2263 -770 -2253
rect -746 -2263 -742 -2253
rect -738 -2263 -734 -2253
rect -730 -2263 -726 -2253
rect -702 -2263 -698 -2253
rect -694 -2263 -690 -2253
rect -686 -2263 -682 -2253
rect -651 -2263 -647 -2253
rect -643 -2263 -639 -2253
rect -287 -2421 -283 -2415
rect -279 -2421 -275 -2415
rect -248 -2470 -244 -2458
rect -230 -2470 -226 -2458
rect -220 -2470 -216 -2458
rect -202 -2470 -198 -2458
rect 3644 -2463 3648 -2457
rect 3652 -2463 3656 -2457
rect -287 -2476 -283 -2470
rect -279 -2476 -275 -2470
rect -754 -2498 -750 -2488
rect -746 -2498 -742 -2488
rect -718 -2498 -714 -2488
rect -710 -2498 -706 -2488
rect -702 -2498 -698 -2488
rect -674 -2498 -670 -2488
rect -666 -2498 -662 -2488
rect -658 -2498 -654 -2488
rect -623 -2498 -619 -2488
rect -615 -2498 -611 -2488
rect 4060 -2483 4064 -2473
rect 4068 -2483 4072 -2473
rect 4096 -2483 4100 -2473
rect 4104 -2483 4108 -2473
rect 4112 -2483 4116 -2473
rect 4140 -2483 4144 -2473
rect 4148 -2483 4152 -2473
rect 4156 -2483 4160 -2473
rect 4191 -2483 4195 -2473
rect 4199 -2483 4203 -2473
rect 3683 -2512 3687 -2500
rect 3701 -2512 3705 -2500
rect 3711 -2512 3715 -2500
rect 3729 -2512 3733 -2500
rect 3644 -2518 3648 -2512
rect 3652 -2518 3656 -2512
rect 187 -2611 191 -2591
rect 206 -2611 210 -2591
rect 229 -2593 233 -2583
rect 237 -2593 241 -2583
rect -745 -2623 -741 -2613
rect -737 -2623 -733 -2613
rect -709 -2623 -705 -2613
rect -701 -2623 -697 -2613
rect -693 -2623 -689 -2613
rect -665 -2623 -661 -2613
rect -657 -2623 -653 -2613
rect -649 -2623 -645 -2613
rect -614 -2623 -610 -2613
rect -606 -2623 -602 -2613
rect 4073 -2775 4077 -2765
rect 4081 -2775 4085 -2765
rect 4109 -2775 4113 -2765
rect 4117 -2775 4121 -2765
rect 4125 -2775 4129 -2765
rect 4153 -2775 4157 -2765
rect 4161 -2775 4165 -2765
rect 4169 -2775 4173 -2765
rect 4204 -2775 4208 -2765
rect 4212 -2775 4216 -2765
rect 3601 -2999 3605 -2993
rect 3609 -2999 3613 -2993
rect 3640 -3048 3644 -3036
rect 3658 -3048 3662 -3036
rect 3668 -3048 3672 -3036
rect 3686 -3048 3690 -3036
rect 3601 -3054 3605 -3048
rect 3609 -3054 3613 -3048
rect 4095 -3149 4099 -3139
rect 4103 -3149 4107 -3139
rect 4131 -3149 4135 -3139
rect 4139 -3149 4143 -3139
rect 4147 -3149 4151 -3139
rect 4175 -3149 4179 -3139
rect 4183 -3149 4187 -3139
rect 4191 -3149 4195 -3139
rect 4226 -3149 4230 -3139
rect 4234 -3149 4238 -3139
<< pdcontact >>
rect -827 -994 -823 -969
rect -819 -994 -815 -969
rect -811 -994 -807 -969
rect -789 -994 -785 -969
rect -781 -994 -777 -969
rect -745 -994 -741 -969
rect -737 -994 -733 -969
rect -700 -994 -696 -969
rect -692 -994 -688 -969
rect -833 -1163 -829 -1138
rect -825 -1163 -821 -1138
rect -817 -1163 -813 -1138
rect -795 -1163 -791 -1138
rect -787 -1163 -783 -1138
rect -751 -1163 -747 -1138
rect -743 -1163 -739 -1138
rect -706 -1163 -702 -1138
rect -698 -1163 -694 -1138
rect 3664 -1203 3668 -1191
rect 3672 -1203 3676 -1191
rect 3703 -1219 3707 -1195
rect 3712 -1219 3716 -1195
rect 3721 -1219 3725 -1195
rect 3731 -1225 3735 -1201
rect 3740 -1225 3744 -1201
rect 3749 -1225 3753 -1201
rect 3664 -1258 3668 -1246
rect 3672 -1258 3676 -1246
rect -833 -1343 -829 -1318
rect -825 -1343 -821 -1318
rect -817 -1343 -813 -1318
rect -795 -1343 -791 -1318
rect -787 -1343 -783 -1318
rect -751 -1343 -747 -1318
rect -743 -1343 -739 -1318
rect -706 -1343 -702 -1318
rect -698 -1343 -694 -1318
rect -298 -1340 -294 -1328
rect -290 -1340 -286 -1328
rect -259 -1356 -255 -1332
rect -250 -1356 -246 -1332
rect -241 -1356 -237 -1332
rect -231 -1362 -227 -1338
rect -222 -1362 -218 -1338
rect -213 -1362 -209 -1338
rect -298 -1395 -294 -1383
rect -290 -1395 -286 -1383
rect 1400 -1476 1404 -1426
rect 1408 -1476 1412 -1426
rect 1450 -1475 1454 -1425
rect 1458 -1475 1462 -1425
rect 1500 -1475 1504 -1425
rect 1508 -1475 1512 -1425
rect 1547 -1475 1551 -1425
rect 1555 -1475 1559 -1425
rect 4094 -1457 4098 -1432
rect 4102 -1457 4106 -1432
rect 4110 -1457 4114 -1432
rect 4132 -1457 4136 -1432
rect 4140 -1457 4144 -1432
rect 4176 -1457 4180 -1432
rect 4184 -1457 4188 -1432
rect 4221 -1457 4225 -1432
rect 4229 -1457 4233 -1432
rect 189 -1554 193 -1534
rect 200 -1554 204 -1534
rect 208 -1554 212 -1534
rect 231 -1561 235 -1541
rect 239 -1561 243 -1541
rect -785 -1659 -781 -1634
rect -777 -1659 -773 -1634
rect -769 -1659 -765 -1634
rect -747 -1659 -743 -1634
rect -739 -1659 -735 -1634
rect -703 -1659 -699 -1634
rect -695 -1659 -691 -1634
rect -658 -1659 -654 -1634
rect -650 -1659 -646 -1634
rect -307 -1699 -303 -1687
rect -299 -1699 -295 -1687
rect -268 -1715 -264 -1691
rect -259 -1715 -255 -1691
rect -250 -1715 -246 -1691
rect -240 -1721 -236 -1697
rect -231 -1721 -227 -1697
rect -222 -1721 -218 -1697
rect -307 -1754 -303 -1742
rect -299 -1754 -295 -1742
rect 1869 -1697 1873 -1657
rect 1877 -1697 1881 -1657
rect 1907 -1697 1911 -1657
rect 1915 -1697 1919 -1657
rect 1951 -1697 1955 -1657
rect 1959 -1697 1963 -1657
rect 1989 -1697 1993 -1657
rect 1997 -1697 2001 -1657
rect 2035 -1695 2039 -1655
rect 2043 -1695 2047 -1655
rect -781 -1821 -777 -1796
rect -773 -1821 -769 -1796
rect -765 -1821 -761 -1796
rect -743 -1821 -739 -1796
rect -735 -1821 -731 -1796
rect -699 -1821 -695 -1796
rect -691 -1821 -687 -1796
rect -654 -1821 -650 -1796
rect -646 -1821 -642 -1796
rect 191 -1904 195 -1884
rect 202 -1904 206 -1884
rect 210 -1904 214 -1884
rect 233 -1911 237 -1891
rect 241 -1911 245 -1891
rect 4079 -1898 4083 -1873
rect 4087 -1898 4091 -1873
rect 4095 -1898 4099 -1873
rect 4117 -1898 4121 -1873
rect 4125 -1898 4129 -1873
rect 4161 -1898 4165 -1873
rect 4169 -1898 4173 -1873
rect 4206 -1898 4210 -1873
rect 4214 -1898 4218 -1873
rect 3704 -2013 3708 -2001
rect 3712 -2013 3716 -2001
rect 3743 -2029 3747 -2005
rect 3752 -2029 3756 -2005
rect 3761 -2029 3765 -2005
rect 3771 -2035 3775 -2011
rect 3780 -2035 3784 -2011
rect 3789 -2035 3793 -2011
rect -776 -2071 -772 -2046
rect -768 -2071 -764 -2046
rect -760 -2071 -756 -2046
rect -738 -2071 -734 -2046
rect -730 -2071 -726 -2046
rect -694 -2071 -690 -2046
rect -686 -2071 -682 -2046
rect -649 -2071 -645 -2046
rect -641 -2071 -637 -2046
rect -280 -2058 -276 -2046
rect -272 -2058 -268 -2046
rect -241 -2074 -237 -2050
rect -232 -2074 -228 -2050
rect -223 -2074 -219 -2050
rect -213 -2080 -209 -2056
rect -204 -2080 -200 -2056
rect -195 -2080 -191 -2056
rect 3704 -2068 3708 -2056
rect 3712 -2068 3716 -2056
rect -280 -2113 -276 -2101
rect -272 -2113 -268 -2101
rect 199 -2196 203 -2176
rect 210 -2196 214 -2176
rect 218 -2196 222 -2176
rect -778 -2231 -774 -2206
rect -770 -2231 -766 -2206
rect -762 -2231 -758 -2206
rect -740 -2231 -736 -2206
rect -732 -2231 -728 -2206
rect -696 -2231 -692 -2206
rect -688 -2231 -684 -2206
rect -651 -2231 -647 -2206
rect -643 -2231 -639 -2206
rect 241 -2203 245 -2183
rect 249 -2203 253 -2183
rect -287 -2401 -283 -2389
rect -279 -2401 -275 -2389
rect -248 -2417 -244 -2393
rect -239 -2417 -235 -2393
rect -230 -2417 -226 -2393
rect -220 -2423 -216 -2399
rect -211 -2423 -207 -2399
rect -202 -2423 -198 -2399
rect -750 -2466 -746 -2441
rect -742 -2466 -738 -2441
rect -734 -2466 -730 -2441
rect -712 -2466 -708 -2441
rect -704 -2466 -700 -2441
rect -668 -2466 -664 -2441
rect -660 -2466 -656 -2441
rect -623 -2466 -619 -2441
rect -615 -2466 -611 -2441
rect -287 -2456 -283 -2444
rect -279 -2456 -275 -2444
rect 3644 -2443 3648 -2431
rect 3652 -2443 3656 -2431
rect 3683 -2459 3687 -2435
rect 3692 -2459 3696 -2435
rect 3701 -2459 3705 -2435
rect 3711 -2465 3715 -2441
rect 3720 -2465 3724 -2441
rect 3729 -2465 3733 -2441
rect 4064 -2451 4068 -2426
rect 4072 -2451 4076 -2426
rect 4080 -2451 4084 -2426
rect 4102 -2451 4106 -2426
rect 4110 -2451 4114 -2426
rect 4146 -2451 4150 -2426
rect 4154 -2451 4158 -2426
rect 4191 -2451 4195 -2426
rect 4199 -2451 4203 -2426
rect 3644 -2498 3648 -2486
rect 3652 -2498 3656 -2486
rect 187 -2562 191 -2542
rect 198 -2562 202 -2542
rect 206 -2562 210 -2542
rect -741 -2591 -737 -2566
rect -733 -2591 -729 -2566
rect -725 -2591 -721 -2566
rect -703 -2591 -699 -2566
rect -695 -2591 -691 -2566
rect -659 -2591 -655 -2566
rect -651 -2591 -647 -2566
rect -614 -2591 -610 -2566
rect -606 -2591 -602 -2566
rect 229 -2569 233 -2549
rect 237 -2569 241 -2549
rect 4077 -2743 4081 -2718
rect 4085 -2743 4089 -2718
rect 4093 -2743 4097 -2718
rect 4115 -2743 4119 -2718
rect 4123 -2743 4127 -2718
rect 4159 -2743 4163 -2718
rect 4167 -2743 4171 -2718
rect 4204 -2743 4208 -2718
rect 4212 -2743 4216 -2718
rect 3601 -2979 3605 -2967
rect 3609 -2979 3613 -2967
rect 3640 -2995 3644 -2971
rect 3649 -2995 3653 -2971
rect 3658 -2995 3662 -2971
rect 3668 -3001 3672 -2977
rect 3677 -3001 3681 -2977
rect 3686 -3001 3690 -2977
rect 3601 -3034 3605 -3022
rect 3609 -3034 3613 -3022
rect 4099 -3117 4103 -3092
rect 4107 -3117 4111 -3092
rect 4115 -3117 4119 -3092
rect 4137 -3117 4141 -3092
rect 4145 -3117 4149 -3092
rect 4181 -3117 4185 -3092
rect 4189 -3117 4193 -3092
rect 4226 -3117 4230 -3092
rect 4234 -3117 4238 -3092
<< psubstratepcontact >>
rect 245 -1594 250 -1590
rect 247 -1944 252 -1940
rect 255 -2236 260 -2232
rect 243 -2602 248 -2598
<< nsubstratencontact >>
rect 1395 -1420 1399 -1415
rect 1445 -1419 1449 -1414
rect 1495 -1419 1499 -1414
rect 1542 -1419 1546 -1414
rect 189 -1529 193 -1523
rect 241 -1534 245 -1530
rect 1864 -1651 1868 -1647
rect 1902 -1651 1906 -1647
rect 1946 -1651 1950 -1647
rect 1984 -1651 1988 -1647
rect 2030 -1649 2034 -1645
rect 191 -1879 195 -1873
rect 243 -1884 247 -1880
rect 199 -2171 203 -2165
rect 251 -2176 255 -2172
rect 187 -2537 191 -2531
rect 239 -2542 243 -2538
<< polysilicon >>
rect -822 -969 -820 -966
rect -814 -969 -812 -966
rect -784 -969 -782 -966
rect -740 -969 -738 -966
rect -695 -969 -693 -966
rect -822 -1001 -820 -994
rect -827 -1005 -820 -1001
rect -826 -1016 -824 -1005
rect -814 -1013 -812 -994
rect -784 -1002 -782 -994
rect -740 -1002 -738 -994
rect -790 -1004 -782 -1002
rect -746 -1004 -738 -1002
rect -790 -1016 -788 -1004
rect -782 -1016 -780 -1007
rect -746 -1016 -744 -1004
rect -738 -1016 -736 -1007
rect -695 -1016 -693 -994
rect -826 -1029 -824 -1026
rect -790 -1029 -788 -1026
rect -782 -1029 -780 -1026
rect -746 -1029 -744 -1026
rect -738 -1029 -736 -1026
rect -695 -1029 -693 -1026
rect -828 -1138 -826 -1135
rect -820 -1138 -818 -1135
rect -790 -1138 -788 -1135
rect -746 -1138 -744 -1135
rect -701 -1138 -699 -1135
rect -828 -1170 -826 -1163
rect -833 -1174 -826 -1170
rect -832 -1185 -830 -1174
rect -820 -1182 -818 -1163
rect -790 -1171 -788 -1163
rect -746 -1171 -744 -1163
rect -796 -1173 -788 -1171
rect -752 -1173 -744 -1171
rect -796 -1185 -794 -1173
rect -788 -1185 -786 -1176
rect -752 -1185 -750 -1173
rect -744 -1185 -742 -1176
rect -701 -1185 -699 -1163
rect 3669 -1191 3671 -1188
rect -832 -1198 -830 -1195
rect -796 -1198 -794 -1195
rect -788 -1198 -786 -1195
rect -752 -1198 -750 -1195
rect -744 -1198 -742 -1195
rect -701 -1198 -699 -1195
rect 3708 -1195 3710 -1192
rect 3718 -1195 3720 -1192
rect 3669 -1217 3671 -1203
rect 3736 -1201 3738 -1198
rect 3746 -1201 3748 -1198
rect 3669 -1226 3671 -1223
rect 3708 -1228 3710 -1219
rect 3718 -1229 3720 -1219
rect 3669 -1246 3671 -1243
rect 3669 -1272 3671 -1258
rect 3708 -1260 3710 -1233
rect 3718 -1260 3720 -1234
rect 3736 -1236 3738 -1225
rect 3736 -1260 3738 -1240
rect 3746 -1247 3748 -1225
rect 3746 -1260 3748 -1251
rect 3708 -1275 3710 -1272
rect 3718 -1275 3720 -1272
rect 3736 -1275 3738 -1272
rect 3746 -1275 3748 -1272
rect 3669 -1281 3671 -1278
rect -828 -1318 -826 -1315
rect -820 -1318 -818 -1315
rect -790 -1318 -788 -1315
rect -746 -1318 -744 -1315
rect -701 -1318 -699 -1315
rect -293 -1328 -291 -1325
rect -254 -1332 -252 -1329
rect -244 -1332 -242 -1329
rect -828 -1350 -826 -1343
rect -833 -1354 -826 -1350
rect -832 -1365 -830 -1354
rect -820 -1362 -818 -1343
rect -790 -1351 -788 -1343
rect -746 -1351 -744 -1343
rect -796 -1353 -788 -1351
rect -752 -1353 -744 -1351
rect -796 -1365 -794 -1353
rect -788 -1365 -786 -1356
rect -752 -1365 -750 -1353
rect -744 -1365 -742 -1356
rect -701 -1365 -699 -1343
rect -293 -1354 -291 -1340
rect -226 -1338 -224 -1335
rect -216 -1338 -214 -1335
rect -293 -1363 -291 -1360
rect -254 -1365 -252 -1356
rect -244 -1366 -242 -1356
rect -832 -1378 -830 -1375
rect -796 -1378 -794 -1375
rect -788 -1378 -786 -1375
rect -752 -1378 -750 -1375
rect -744 -1378 -742 -1375
rect -701 -1378 -699 -1375
rect -293 -1383 -291 -1380
rect -293 -1409 -291 -1395
rect -254 -1397 -252 -1370
rect -244 -1397 -242 -1371
rect -226 -1373 -224 -1362
rect -226 -1397 -224 -1377
rect -216 -1384 -214 -1362
rect -216 -1397 -214 -1388
rect -254 -1412 -252 -1409
rect -244 -1412 -242 -1409
rect -226 -1412 -224 -1409
rect -216 -1412 -214 -1409
rect -293 -1418 -291 -1415
rect 1405 -1426 1407 -1423
rect 1455 -1425 1457 -1422
rect 1505 -1425 1507 -1422
rect 1552 -1425 1554 -1422
rect 4099 -1432 4101 -1429
rect 4107 -1432 4109 -1429
rect 4137 -1432 4139 -1429
rect 4181 -1432 4183 -1429
rect 4226 -1432 4228 -1429
rect 4099 -1464 4101 -1457
rect 4094 -1468 4101 -1464
rect 1405 -1499 1407 -1476
rect 1455 -1498 1457 -1475
rect 1505 -1498 1507 -1475
rect 1552 -1498 1554 -1475
rect 4095 -1479 4097 -1468
rect 4107 -1476 4109 -1457
rect 4137 -1465 4139 -1457
rect 4181 -1465 4183 -1457
rect 4131 -1467 4139 -1465
rect 4175 -1467 4183 -1465
rect 4131 -1479 4133 -1467
rect 4139 -1479 4141 -1470
rect 4175 -1479 4177 -1467
rect 4183 -1479 4185 -1470
rect 4226 -1479 4228 -1457
rect 4095 -1492 4097 -1489
rect 4131 -1492 4133 -1489
rect 4139 -1492 4141 -1489
rect 4175 -1492 4177 -1489
rect 4183 -1492 4185 -1489
rect 4226 -1492 4228 -1489
rect 194 -1534 196 -1531
rect 205 -1534 207 -1531
rect 236 -1541 238 -1537
rect 194 -1583 196 -1554
rect 205 -1583 207 -1554
rect 236 -1575 238 -1561
rect 236 -1588 238 -1585
rect 194 -1606 196 -1603
rect 205 -1606 207 -1603
rect -780 -1634 -778 -1631
rect -772 -1634 -770 -1631
rect -742 -1634 -740 -1631
rect -698 -1634 -696 -1631
rect -653 -1634 -651 -1631
rect 1874 -1657 1876 -1654
rect 1912 -1657 1914 -1654
rect 1956 -1657 1958 -1654
rect 1994 -1657 1996 -1654
rect 2040 -1655 2042 -1652
rect -780 -1666 -778 -1659
rect -785 -1670 -778 -1666
rect -784 -1681 -782 -1670
rect -772 -1678 -770 -1659
rect -742 -1667 -740 -1659
rect -698 -1667 -696 -1659
rect -748 -1669 -740 -1667
rect -704 -1669 -696 -1667
rect -748 -1681 -746 -1669
rect -740 -1681 -738 -1672
rect -704 -1681 -702 -1669
rect -696 -1681 -694 -1672
rect -653 -1681 -651 -1659
rect 1341 -1662 1343 -1659
rect 1369 -1662 1371 -1659
rect 1396 -1662 1398 -1659
rect 1435 -1662 1437 -1659
rect 1463 -1662 1465 -1659
rect 1490 -1662 1492 -1659
rect 1530 -1661 1532 -1658
rect 1558 -1661 1560 -1658
rect 1585 -1661 1587 -1658
rect 1621 -1661 1623 -1658
rect -302 -1687 -300 -1684
rect -784 -1694 -782 -1691
rect -748 -1694 -746 -1691
rect -740 -1694 -738 -1691
rect -704 -1694 -702 -1691
rect -696 -1694 -694 -1691
rect -653 -1694 -651 -1691
rect -263 -1691 -261 -1688
rect -253 -1691 -251 -1688
rect -302 -1713 -300 -1699
rect -235 -1697 -233 -1694
rect -225 -1697 -223 -1694
rect -302 -1722 -300 -1719
rect -263 -1724 -261 -1715
rect -253 -1725 -251 -1715
rect -302 -1742 -300 -1739
rect -302 -1768 -300 -1754
rect -263 -1756 -261 -1729
rect -253 -1756 -251 -1730
rect -235 -1732 -233 -1721
rect -235 -1756 -233 -1736
rect -225 -1743 -223 -1721
rect -225 -1756 -223 -1747
rect 1874 -1715 1876 -1697
rect 1912 -1715 1914 -1697
rect 1956 -1715 1958 -1697
rect 1994 -1715 1996 -1697
rect 2040 -1713 2042 -1695
rect 1874 -1739 1876 -1735
rect 1912 -1739 1914 -1735
rect 1956 -1739 1958 -1735
rect 1994 -1739 1996 -1735
rect 2040 -1737 2042 -1733
rect -263 -1771 -261 -1768
rect -253 -1771 -251 -1768
rect -235 -1771 -233 -1768
rect -225 -1771 -223 -1768
rect 1341 -1774 1343 -1762
rect 1369 -1774 1371 -1762
rect 1396 -1774 1398 -1762
rect 1435 -1774 1437 -1762
rect 1463 -1774 1465 -1762
rect 1490 -1774 1492 -1762
rect 1530 -1773 1532 -1761
rect 1558 -1773 1560 -1761
rect 1585 -1773 1587 -1761
rect 1621 -1773 1623 -1761
rect -302 -1777 -300 -1774
rect -776 -1796 -774 -1793
rect -768 -1796 -766 -1793
rect -738 -1796 -736 -1793
rect -694 -1796 -692 -1793
rect -649 -1796 -647 -1793
rect -776 -1828 -774 -1821
rect -781 -1832 -774 -1828
rect -780 -1843 -778 -1832
rect -768 -1840 -766 -1821
rect -738 -1829 -736 -1821
rect -694 -1829 -692 -1821
rect -744 -1831 -736 -1829
rect -700 -1831 -692 -1829
rect -744 -1843 -742 -1831
rect -736 -1843 -734 -1834
rect -700 -1843 -698 -1831
rect -692 -1843 -690 -1834
rect -649 -1843 -647 -1821
rect -780 -1856 -778 -1853
rect -744 -1856 -742 -1853
rect -736 -1856 -734 -1853
rect -700 -1856 -698 -1853
rect -692 -1856 -690 -1853
rect -649 -1856 -647 -1853
rect 4084 -1873 4086 -1870
rect 4092 -1873 4094 -1870
rect 4122 -1873 4124 -1870
rect 4166 -1873 4168 -1870
rect 4211 -1873 4213 -1870
rect 196 -1884 198 -1881
rect 207 -1884 209 -1881
rect 238 -1891 240 -1887
rect 196 -1933 198 -1904
rect 207 -1933 209 -1904
rect 4084 -1905 4086 -1898
rect 4079 -1909 4086 -1905
rect 238 -1925 240 -1911
rect 4080 -1920 4082 -1909
rect 4092 -1917 4094 -1898
rect 4122 -1906 4124 -1898
rect 4166 -1906 4168 -1898
rect 4116 -1908 4124 -1906
rect 4160 -1908 4168 -1906
rect 4116 -1920 4118 -1908
rect 4124 -1920 4126 -1911
rect 4160 -1920 4162 -1908
rect 4168 -1920 4170 -1911
rect 4211 -1920 4213 -1898
rect 4080 -1933 4082 -1930
rect 4116 -1933 4118 -1930
rect 4124 -1933 4126 -1930
rect 4160 -1933 4162 -1930
rect 4168 -1933 4170 -1930
rect 4211 -1933 4213 -1930
rect 238 -1938 240 -1935
rect 196 -1956 198 -1953
rect 207 -1956 209 -1953
rect 3709 -2001 3711 -1998
rect 3748 -2005 3750 -2002
rect 3758 -2005 3760 -2002
rect 3709 -2027 3711 -2013
rect 3776 -2011 3778 -2008
rect 3786 -2011 3788 -2008
rect 3709 -2036 3711 -2033
rect 3748 -2038 3750 -2029
rect 3758 -2039 3760 -2029
rect -771 -2046 -769 -2043
rect -763 -2046 -761 -2043
rect -733 -2046 -731 -2043
rect -689 -2046 -687 -2043
rect -644 -2046 -642 -2043
rect -275 -2046 -273 -2043
rect -236 -2050 -234 -2047
rect -226 -2050 -224 -2047
rect -771 -2078 -769 -2071
rect -776 -2082 -769 -2078
rect -775 -2093 -773 -2082
rect -763 -2090 -761 -2071
rect -733 -2079 -731 -2071
rect -689 -2079 -687 -2071
rect -739 -2081 -731 -2079
rect -695 -2081 -687 -2079
rect -739 -2093 -737 -2081
rect -731 -2093 -729 -2084
rect -695 -2093 -693 -2081
rect -687 -2093 -685 -2084
rect -644 -2093 -642 -2071
rect -275 -2072 -273 -2058
rect -208 -2056 -206 -2053
rect -198 -2056 -196 -2053
rect 3709 -2056 3711 -2053
rect -275 -2081 -273 -2078
rect -236 -2083 -234 -2074
rect -226 -2084 -224 -2074
rect -275 -2101 -273 -2098
rect -775 -2106 -773 -2103
rect -739 -2106 -737 -2103
rect -731 -2106 -729 -2103
rect -695 -2106 -693 -2103
rect -687 -2106 -685 -2103
rect -644 -2106 -642 -2103
rect -275 -2127 -273 -2113
rect -236 -2115 -234 -2088
rect -226 -2115 -224 -2089
rect -208 -2091 -206 -2080
rect -208 -2115 -206 -2095
rect -198 -2102 -196 -2080
rect 3709 -2082 3711 -2068
rect 3748 -2070 3750 -2043
rect 3758 -2070 3760 -2044
rect 3776 -2046 3778 -2035
rect 3776 -2070 3778 -2050
rect 3786 -2057 3788 -2035
rect 3786 -2070 3788 -2061
rect 3748 -2085 3750 -2082
rect 3758 -2085 3760 -2082
rect 3776 -2085 3778 -2082
rect 3786 -2085 3788 -2082
rect 3709 -2091 3711 -2088
rect -198 -2115 -196 -2106
rect -236 -2130 -234 -2127
rect -226 -2130 -224 -2127
rect -208 -2130 -206 -2127
rect -198 -2130 -196 -2127
rect -275 -2136 -273 -2133
rect 204 -2176 206 -2173
rect 215 -2176 217 -2173
rect 246 -2183 248 -2179
rect -773 -2206 -771 -2203
rect -765 -2206 -763 -2203
rect -735 -2206 -733 -2203
rect -691 -2206 -689 -2203
rect -646 -2206 -644 -2203
rect 204 -2225 206 -2196
rect 215 -2225 217 -2196
rect 246 -2217 248 -2203
rect -773 -2238 -771 -2231
rect -778 -2242 -771 -2238
rect -777 -2253 -775 -2242
rect -765 -2250 -763 -2231
rect -735 -2239 -733 -2231
rect -691 -2239 -689 -2231
rect -741 -2241 -733 -2239
rect -697 -2241 -689 -2239
rect -741 -2253 -739 -2241
rect -733 -2253 -731 -2244
rect -697 -2253 -695 -2241
rect -689 -2253 -687 -2244
rect -646 -2253 -644 -2231
rect 246 -2230 248 -2227
rect 204 -2248 206 -2245
rect 215 -2248 217 -2245
rect -777 -2266 -775 -2263
rect -741 -2266 -739 -2263
rect -733 -2266 -731 -2263
rect -697 -2266 -695 -2263
rect -689 -2266 -687 -2263
rect -646 -2266 -644 -2263
rect -282 -2389 -280 -2386
rect -243 -2393 -241 -2390
rect -233 -2393 -231 -2390
rect -282 -2415 -280 -2401
rect -215 -2399 -213 -2396
rect -205 -2399 -203 -2396
rect -282 -2424 -280 -2421
rect -243 -2426 -241 -2417
rect -233 -2427 -231 -2417
rect -745 -2441 -743 -2438
rect -737 -2441 -735 -2438
rect -707 -2441 -705 -2438
rect -663 -2441 -661 -2438
rect -618 -2441 -616 -2438
rect -282 -2444 -280 -2441
rect -745 -2473 -743 -2466
rect -750 -2477 -743 -2473
rect -749 -2488 -747 -2477
rect -737 -2485 -735 -2466
rect -707 -2474 -705 -2466
rect -663 -2474 -661 -2466
rect -713 -2476 -705 -2474
rect -669 -2476 -661 -2474
rect -713 -2488 -711 -2476
rect -705 -2488 -703 -2479
rect -669 -2488 -667 -2476
rect -661 -2488 -659 -2479
rect -618 -2488 -616 -2466
rect -282 -2470 -280 -2456
rect -243 -2458 -241 -2431
rect -233 -2458 -231 -2432
rect -215 -2434 -213 -2423
rect -215 -2458 -213 -2438
rect -205 -2445 -203 -2423
rect 4069 -2426 4071 -2423
rect 4077 -2426 4079 -2423
rect 4107 -2426 4109 -2423
rect 4151 -2426 4153 -2423
rect 4196 -2426 4198 -2423
rect 3649 -2431 3651 -2428
rect 3688 -2435 3690 -2432
rect 3698 -2435 3700 -2432
rect -205 -2458 -203 -2449
rect 3649 -2457 3651 -2443
rect 3716 -2441 3718 -2438
rect 3726 -2441 3728 -2438
rect 3649 -2466 3651 -2463
rect 3688 -2468 3690 -2459
rect -243 -2473 -241 -2470
rect -233 -2473 -231 -2470
rect -215 -2473 -213 -2470
rect -205 -2473 -203 -2470
rect 3698 -2469 3700 -2459
rect 4069 -2458 4071 -2451
rect 4064 -2462 4071 -2458
rect -282 -2479 -280 -2476
rect 3649 -2486 3651 -2483
rect -749 -2501 -747 -2498
rect -713 -2501 -711 -2498
rect -705 -2501 -703 -2498
rect -669 -2501 -667 -2498
rect -661 -2501 -659 -2498
rect -618 -2501 -616 -2498
rect 3649 -2512 3651 -2498
rect 3688 -2500 3690 -2473
rect 3698 -2500 3700 -2474
rect 3716 -2476 3718 -2465
rect 3716 -2500 3718 -2480
rect 3726 -2487 3728 -2465
rect 4065 -2473 4067 -2462
rect 4077 -2470 4079 -2451
rect 4107 -2459 4109 -2451
rect 4151 -2459 4153 -2451
rect 4101 -2461 4109 -2459
rect 4145 -2461 4153 -2459
rect 4101 -2473 4103 -2461
rect 4109 -2473 4111 -2464
rect 4145 -2473 4147 -2461
rect 4153 -2473 4155 -2464
rect 4196 -2473 4198 -2451
rect 4065 -2486 4067 -2483
rect 4101 -2486 4103 -2483
rect 4109 -2486 4111 -2483
rect 4145 -2486 4147 -2483
rect 4153 -2486 4155 -2483
rect 4196 -2486 4198 -2483
rect 3726 -2500 3728 -2491
rect 3688 -2515 3690 -2512
rect 3698 -2515 3700 -2512
rect 3716 -2515 3718 -2512
rect 3726 -2515 3728 -2512
rect 3649 -2521 3651 -2518
rect 192 -2542 194 -2539
rect 203 -2542 205 -2539
rect 234 -2549 236 -2545
rect -736 -2566 -734 -2563
rect -728 -2566 -726 -2563
rect -698 -2566 -696 -2563
rect -654 -2566 -652 -2563
rect -609 -2566 -607 -2563
rect 192 -2591 194 -2562
rect 203 -2591 205 -2562
rect 234 -2583 236 -2569
rect -736 -2598 -734 -2591
rect -741 -2602 -734 -2598
rect -740 -2613 -738 -2602
rect -728 -2610 -726 -2591
rect -698 -2599 -696 -2591
rect -654 -2599 -652 -2591
rect -704 -2601 -696 -2599
rect -660 -2601 -652 -2599
rect -704 -2613 -702 -2601
rect -696 -2613 -694 -2604
rect -660 -2613 -658 -2601
rect -652 -2613 -650 -2604
rect -609 -2613 -607 -2591
rect 234 -2596 236 -2593
rect 192 -2614 194 -2611
rect 203 -2614 205 -2611
rect -740 -2626 -738 -2623
rect -704 -2626 -702 -2623
rect -696 -2626 -694 -2623
rect -660 -2626 -658 -2623
rect -652 -2626 -650 -2623
rect -609 -2626 -607 -2623
rect 4082 -2718 4084 -2715
rect 4090 -2718 4092 -2715
rect 4120 -2718 4122 -2715
rect 4164 -2718 4166 -2715
rect 4209 -2718 4211 -2715
rect 4082 -2750 4084 -2743
rect 4077 -2754 4084 -2750
rect 4078 -2765 4080 -2754
rect 4090 -2762 4092 -2743
rect 4120 -2751 4122 -2743
rect 4164 -2751 4166 -2743
rect 4114 -2753 4122 -2751
rect 4158 -2753 4166 -2751
rect 4114 -2765 4116 -2753
rect 4122 -2765 4124 -2756
rect 4158 -2765 4160 -2753
rect 4166 -2765 4168 -2756
rect 4209 -2765 4211 -2743
rect 4078 -2778 4080 -2775
rect 4114 -2778 4116 -2775
rect 4122 -2778 4124 -2775
rect 4158 -2778 4160 -2775
rect 4166 -2778 4168 -2775
rect 4209 -2778 4211 -2775
rect 3606 -2967 3608 -2964
rect 3645 -2971 3647 -2968
rect 3655 -2971 3657 -2968
rect 3606 -2993 3608 -2979
rect 3673 -2977 3675 -2974
rect 3683 -2977 3685 -2974
rect 3606 -3002 3608 -2999
rect 3645 -3004 3647 -2995
rect 3655 -3005 3657 -2995
rect 3606 -3022 3608 -3019
rect 3606 -3048 3608 -3034
rect 3645 -3036 3647 -3009
rect 3655 -3036 3657 -3010
rect 3673 -3012 3675 -3001
rect 3673 -3036 3675 -3016
rect 3683 -3023 3685 -3001
rect 3683 -3036 3685 -3027
rect 3645 -3051 3647 -3048
rect 3655 -3051 3657 -3048
rect 3673 -3051 3675 -3048
rect 3683 -3051 3685 -3048
rect 3606 -3057 3608 -3054
rect 4104 -3092 4106 -3089
rect 4112 -3092 4114 -3089
rect 4142 -3092 4144 -3089
rect 4186 -3092 4188 -3089
rect 4231 -3092 4233 -3089
rect 4104 -3124 4106 -3117
rect 4099 -3128 4106 -3124
rect 4100 -3139 4102 -3128
rect 4112 -3136 4114 -3117
rect 4142 -3125 4144 -3117
rect 4186 -3125 4188 -3117
rect 4136 -3127 4144 -3125
rect 4180 -3127 4188 -3125
rect 4136 -3139 4138 -3127
rect 4144 -3139 4146 -3130
rect 4180 -3139 4182 -3127
rect 4188 -3139 4190 -3130
rect 4231 -3139 4233 -3117
rect 4100 -3152 4102 -3149
rect 4136 -3152 4138 -3149
rect 4144 -3152 4146 -3149
rect 4180 -3152 4182 -3149
rect 4188 -3152 4190 -3149
rect 4231 -3152 4233 -3149
<< polycontact >>
rect -831 -1005 -827 -1001
rect -818 -1013 -814 -1009
rect -807 -1005 -803 -1001
rect -795 -1013 -790 -1008
rect -780 -1013 -776 -1009
rect -751 -1013 -746 -1008
rect -699 -1008 -695 -1003
rect -736 -1013 -732 -1009
rect -837 -1174 -833 -1170
rect -824 -1182 -820 -1178
rect -813 -1174 -809 -1170
rect -801 -1182 -796 -1177
rect -786 -1182 -782 -1178
rect -757 -1182 -752 -1177
rect -705 -1177 -701 -1172
rect -742 -1182 -738 -1178
rect 3665 -1214 3669 -1210
rect 3665 -1269 3669 -1265
rect 3734 -1240 3738 -1236
rect 3745 -1251 3749 -1247
rect -837 -1354 -833 -1350
rect -824 -1362 -820 -1358
rect -813 -1354 -809 -1350
rect -801 -1362 -796 -1357
rect -786 -1362 -782 -1358
rect -757 -1362 -752 -1357
rect -705 -1357 -701 -1352
rect -742 -1362 -738 -1358
rect -297 -1351 -293 -1347
rect -297 -1406 -293 -1402
rect -228 -1377 -224 -1373
rect -217 -1388 -213 -1384
rect 4090 -1468 4094 -1464
rect 4103 -1476 4107 -1472
rect 4114 -1468 4118 -1464
rect 4126 -1476 4131 -1471
rect 4141 -1476 4145 -1472
rect 4170 -1476 4175 -1471
rect 4222 -1471 4226 -1466
rect 4185 -1476 4189 -1472
rect 190 -1580 194 -1576
rect 201 -1573 205 -1569
rect 232 -1572 236 -1568
rect -789 -1670 -785 -1666
rect -776 -1678 -772 -1674
rect -765 -1670 -761 -1666
rect -753 -1678 -748 -1673
rect -738 -1678 -734 -1674
rect -709 -1678 -704 -1673
rect -657 -1673 -653 -1668
rect -694 -1678 -690 -1674
rect -306 -1710 -302 -1706
rect -306 -1765 -302 -1761
rect -237 -1736 -233 -1732
rect -226 -1747 -222 -1743
rect -785 -1832 -781 -1828
rect -772 -1840 -768 -1836
rect -761 -1832 -757 -1828
rect -749 -1840 -744 -1835
rect -734 -1840 -730 -1836
rect -705 -1840 -700 -1835
rect -653 -1835 -649 -1830
rect -690 -1840 -686 -1836
rect 192 -1930 196 -1926
rect 203 -1923 207 -1919
rect 4075 -1909 4079 -1905
rect 234 -1922 238 -1918
rect 4088 -1917 4092 -1913
rect 4099 -1909 4103 -1905
rect 4111 -1917 4116 -1912
rect 4126 -1917 4130 -1913
rect 4155 -1917 4160 -1912
rect 4207 -1912 4211 -1907
rect 4170 -1917 4174 -1913
rect 3705 -2024 3709 -2020
rect -279 -2069 -275 -2065
rect -780 -2082 -776 -2078
rect -767 -2090 -763 -2086
rect -756 -2082 -752 -2078
rect -744 -2090 -739 -2085
rect -729 -2090 -725 -2086
rect -700 -2090 -695 -2085
rect -648 -2085 -644 -2080
rect -685 -2090 -681 -2086
rect 3705 -2079 3709 -2075
rect -279 -2124 -275 -2120
rect -210 -2095 -206 -2091
rect 3774 -2050 3778 -2046
rect 3785 -2061 3789 -2057
rect -199 -2106 -195 -2102
rect 200 -2222 204 -2218
rect 211 -2215 215 -2211
rect 242 -2214 246 -2210
rect -782 -2242 -778 -2238
rect -769 -2250 -765 -2246
rect -758 -2242 -754 -2238
rect -746 -2250 -741 -2245
rect -731 -2250 -727 -2246
rect -702 -2250 -697 -2245
rect -650 -2245 -646 -2240
rect -687 -2250 -683 -2246
rect -286 -2412 -282 -2408
rect -754 -2477 -750 -2473
rect -741 -2485 -737 -2481
rect -730 -2477 -726 -2473
rect -718 -2485 -713 -2480
rect -703 -2485 -699 -2481
rect -674 -2485 -669 -2480
rect -622 -2480 -618 -2475
rect -659 -2485 -655 -2481
rect -286 -2467 -282 -2463
rect -217 -2438 -213 -2434
rect -206 -2449 -202 -2445
rect 3645 -2454 3649 -2450
rect 4060 -2462 4064 -2458
rect 3645 -2509 3649 -2505
rect 3714 -2480 3718 -2476
rect 4073 -2470 4077 -2466
rect 4084 -2462 4088 -2458
rect 4096 -2470 4101 -2465
rect 4111 -2470 4115 -2466
rect 4140 -2470 4145 -2465
rect 4192 -2465 4196 -2460
rect 4155 -2470 4159 -2466
rect 3725 -2491 3729 -2487
rect 188 -2588 192 -2584
rect 199 -2581 203 -2577
rect 230 -2580 234 -2576
rect -745 -2602 -741 -2598
rect -732 -2610 -728 -2606
rect -721 -2602 -717 -2598
rect -709 -2610 -704 -2605
rect -694 -2610 -690 -2606
rect -665 -2610 -660 -2605
rect -613 -2605 -609 -2600
rect -650 -2610 -646 -2606
rect 4073 -2754 4077 -2750
rect 4086 -2762 4090 -2758
rect 4097 -2754 4101 -2750
rect 4109 -2762 4114 -2757
rect 4124 -2762 4128 -2758
rect 4153 -2762 4158 -2757
rect 4205 -2757 4209 -2752
rect 4168 -2762 4172 -2758
rect 3602 -2990 3606 -2986
rect 3602 -3045 3606 -3041
rect 3671 -3016 3675 -3012
rect 3682 -3027 3686 -3023
rect 4095 -3128 4099 -3124
rect 4108 -3136 4112 -3132
rect 4119 -3128 4123 -3124
rect 4131 -3136 4136 -3131
rect 4146 -3136 4150 -3132
rect 4175 -3136 4180 -3131
rect 4227 -3131 4231 -3126
rect 4190 -3136 4194 -3132
<< metal1 >>
rect -833 -963 -680 -959
rect -827 -969 -823 -963
rect -789 -969 -785 -963
rect -745 -969 -741 -963
rect -700 -969 -696 -963
rect -777 -994 -764 -969
rect -733 -994 -720 -969
rect -838 -1005 -831 -1001
rect -827 -1013 -818 -1009
rect -811 -1016 -807 -994
rect -803 -1005 -802 -1001
rect -767 -1003 -764 -994
rect -723 -1003 -720 -994
rect -767 -1008 -755 -1003
rect -723 -1008 -699 -1003
rect -692 -1004 -688 -994
rect -803 -1010 -795 -1008
rect -798 -1013 -795 -1010
rect -776 -1013 -775 -1009
rect -767 -1016 -764 -1008
rect -759 -1013 -751 -1008
rect -732 -1013 -731 -1009
rect -723 -1016 -720 -1008
rect -692 -1009 -679 -1004
rect -692 -1016 -688 -1009
rect -819 -1026 -807 -1016
rect -775 -1026 -764 -1016
rect -731 -1026 -720 -1016
rect -831 -1031 -827 -1026
rect -795 -1031 -791 -1026
rect -751 -1031 -747 -1026
rect -700 -1031 -696 -1026
rect -832 -1035 -688 -1031
rect -839 -1132 -686 -1128
rect -833 -1138 -829 -1132
rect -795 -1138 -791 -1132
rect -751 -1138 -747 -1132
rect -706 -1138 -702 -1132
rect -783 -1163 -770 -1138
rect -739 -1163 -726 -1138
rect -844 -1174 -837 -1170
rect -833 -1182 -824 -1178
rect -817 -1185 -813 -1163
rect -809 -1174 -808 -1170
rect -773 -1172 -770 -1163
rect -729 -1172 -726 -1163
rect -773 -1177 -761 -1172
rect -729 -1177 -705 -1172
rect -698 -1173 -694 -1163
rect -809 -1179 -801 -1177
rect -804 -1182 -801 -1179
rect -782 -1182 -781 -1178
rect -773 -1185 -770 -1177
rect -765 -1182 -757 -1177
rect -738 -1182 -737 -1178
rect -729 -1185 -726 -1177
rect -698 -1178 -685 -1173
rect -698 -1185 -694 -1178
rect 3663 -1185 3691 -1182
rect -825 -1195 -813 -1185
rect -781 -1195 -770 -1185
rect -737 -1195 -726 -1185
rect 3664 -1191 3667 -1185
rect 3688 -1186 3691 -1185
rect 3688 -1189 3759 -1186
rect -837 -1200 -833 -1195
rect -801 -1200 -797 -1195
rect -757 -1200 -753 -1195
rect -706 -1200 -702 -1195
rect -838 -1204 -694 -1200
rect 3647 -1215 3650 -1212
rect 3655 -1214 3665 -1211
rect 3673 -1211 3676 -1203
rect 3703 -1195 3706 -1189
rect 3722 -1195 3725 -1189
rect 3673 -1214 3694 -1211
rect 3673 -1217 3676 -1214
rect 3664 -1227 3667 -1223
rect 3658 -1229 3682 -1227
rect 3658 -1230 3676 -1229
rect 3681 -1230 3682 -1229
rect 3691 -1237 3694 -1214
rect 3732 -1195 3752 -1192
rect 3732 -1201 3735 -1195
rect 3749 -1201 3752 -1195
rect 3713 -1222 3716 -1219
rect 3713 -1225 3731 -1222
rect 3741 -1232 3744 -1225
rect 3741 -1235 3758 -1232
rect 3663 -1238 3682 -1237
rect 3658 -1240 3682 -1238
rect 3691 -1240 3734 -1237
rect 3664 -1246 3667 -1240
rect 3755 -1246 3758 -1235
rect 3720 -1251 3745 -1248
rect 3755 -1250 3768 -1246
rect 3720 -1253 3723 -1251
rect 3647 -1269 3650 -1266
rect 3655 -1269 3665 -1266
rect 3673 -1266 3676 -1258
rect 3685 -1256 3723 -1253
rect 3755 -1254 3758 -1250
rect 3685 -1266 3688 -1256
rect 3726 -1257 3758 -1254
rect 3726 -1260 3729 -1257
rect 3673 -1269 3688 -1266
rect 3673 -1272 3676 -1269
rect 3725 -1263 3731 -1260
rect 3664 -1282 3667 -1278
rect 3685 -1279 3690 -1276
rect 3703 -1276 3706 -1272
rect 3750 -1276 3753 -1272
rect 3695 -1279 3759 -1276
rect 3685 -1282 3688 -1279
rect 3658 -1285 3688 -1282
rect 3764 -1290 3768 -1250
rect -839 -1312 -686 -1308
rect -833 -1318 -829 -1312
rect -795 -1318 -791 -1312
rect -751 -1318 -747 -1312
rect -706 -1318 -702 -1312
rect -783 -1343 -770 -1318
rect -739 -1343 -726 -1318
rect -299 -1322 -271 -1319
rect -298 -1328 -295 -1322
rect -274 -1323 -271 -1322
rect -274 -1326 -203 -1323
rect -844 -1354 -837 -1350
rect -833 -1362 -824 -1358
rect -817 -1365 -813 -1343
rect -809 -1354 -808 -1350
rect -773 -1352 -770 -1343
rect -729 -1352 -726 -1343
rect -773 -1357 -761 -1352
rect -729 -1357 -705 -1352
rect -698 -1353 -694 -1343
rect -315 -1352 -312 -1349
rect -307 -1351 -297 -1348
rect -289 -1348 -286 -1340
rect -259 -1332 -256 -1326
rect -240 -1332 -237 -1326
rect -289 -1351 -268 -1348
rect -809 -1359 -801 -1357
rect -804 -1362 -801 -1359
rect -782 -1362 -781 -1358
rect -773 -1365 -770 -1357
rect -765 -1362 -757 -1357
rect -738 -1362 -737 -1358
rect -729 -1365 -726 -1357
rect -698 -1358 -685 -1353
rect -289 -1354 -286 -1351
rect -698 -1365 -694 -1358
rect -298 -1364 -295 -1360
rect -825 -1375 -813 -1365
rect -781 -1375 -770 -1365
rect -737 -1375 -726 -1365
rect -304 -1366 -280 -1364
rect -304 -1367 -286 -1366
rect -281 -1367 -280 -1366
rect -271 -1374 -268 -1351
rect -230 -1332 -210 -1329
rect -230 -1338 -227 -1332
rect -213 -1338 -210 -1332
rect -249 -1359 -246 -1356
rect -249 -1362 -231 -1359
rect -221 -1369 -218 -1362
rect -221 -1372 -204 -1369
rect -299 -1375 -280 -1374
rect -837 -1380 -833 -1375
rect -801 -1380 -797 -1375
rect -757 -1380 -753 -1375
rect -706 -1380 -702 -1375
rect -304 -1377 -280 -1375
rect -271 -1377 -228 -1374
rect -838 -1384 -694 -1380
rect -298 -1383 -295 -1377
rect -207 -1383 -204 -1372
rect -242 -1388 -217 -1385
rect -207 -1387 -194 -1383
rect -242 -1390 -239 -1388
rect -315 -1406 -312 -1403
rect -307 -1406 -297 -1403
rect -289 -1403 -286 -1395
rect -277 -1393 -239 -1390
rect -207 -1391 -204 -1387
rect -277 -1403 -274 -1393
rect -236 -1394 -204 -1391
rect -236 -1397 -233 -1394
rect -289 -1406 -274 -1403
rect -289 -1409 -286 -1406
rect -237 -1400 -231 -1397
rect -298 -1419 -295 -1415
rect -277 -1416 -272 -1413
rect -259 -1413 -256 -1409
rect -212 -1413 -209 -1409
rect -267 -1416 -203 -1413
rect -277 -1419 -274 -1416
rect -304 -1422 -274 -1419
rect -198 -1427 -194 -1387
rect 1400 -1415 1404 -1406
rect 1450 -1414 1454 -1405
rect 1500 -1414 1504 -1405
rect 1547 -1414 1551 -1405
rect 1394 -1420 1395 -1415
rect 1399 -1420 1418 -1415
rect 1444 -1419 1445 -1414
rect 1449 -1419 1468 -1414
rect 1494 -1419 1495 -1414
rect 1499 -1419 1518 -1414
rect 1541 -1419 1542 -1414
rect 1546 -1419 1565 -1414
rect 1400 -1426 1404 -1420
rect 1450 -1425 1454 -1419
rect 1500 -1425 1504 -1419
rect 1547 -1425 1551 -1419
rect 4088 -1426 4241 -1422
rect 4094 -1432 4098 -1426
rect 4132 -1432 4136 -1426
rect 4176 -1432 4180 -1426
rect 4221 -1432 4225 -1426
rect 4144 -1457 4157 -1432
rect 4188 -1457 4201 -1432
rect 4083 -1468 4090 -1464
rect 1408 -1490 1412 -1476
rect 1458 -1489 1462 -1475
rect 1508 -1489 1512 -1475
rect 1555 -1489 1559 -1475
rect 4094 -1476 4103 -1472
rect 4110 -1479 4114 -1457
rect 4118 -1468 4119 -1464
rect 4154 -1466 4157 -1457
rect 4198 -1466 4201 -1457
rect 4154 -1471 4166 -1466
rect 4198 -1471 4222 -1466
rect 4229 -1467 4233 -1457
rect 4118 -1473 4126 -1471
rect 4123 -1476 4126 -1473
rect 4145 -1476 4146 -1472
rect 4154 -1479 4157 -1471
rect 4162 -1476 4170 -1471
rect 4189 -1476 4190 -1472
rect 4198 -1479 4201 -1471
rect 4229 -1472 4242 -1467
rect 4229 -1479 4233 -1472
rect 4102 -1489 4114 -1479
rect 4146 -1489 4157 -1479
rect 4190 -1489 4201 -1479
rect 4090 -1494 4094 -1489
rect 4126 -1494 4130 -1489
rect 4170 -1494 4174 -1489
rect 4221 -1494 4225 -1489
rect 4089 -1498 4233 -1494
rect 189 -1523 212 -1519
rect 193 -1525 212 -1523
rect 189 -1534 193 -1529
rect 208 -1534 212 -1525
rect 225 -1530 249 -1529
rect 225 -1534 241 -1530
rect 245 -1534 249 -1530
rect 225 -1536 249 -1534
rect 231 -1541 235 -1536
rect 200 -1562 204 -1554
rect 200 -1566 212 -1562
rect 208 -1568 212 -1566
rect 239 -1568 243 -1561
rect 183 -1573 201 -1569
rect 208 -1572 232 -1568
rect 239 -1572 249 -1568
rect 183 -1580 190 -1576
rect 208 -1583 212 -1572
rect 239 -1575 243 -1572
rect 231 -1589 235 -1585
rect 225 -1590 250 -1589
rect 225 -1594 245 -1590
rect 225 -1595 250 -1594
rect 189 -1607 193 -1603
rect 189 -1611 205 -1607
rect -791 -1628 -638 -1624
rect -785 -1634 -781 -1628
rect -747 -1634 -743 -1628
rect -703 -1634 -699 -1628
rect -658 -1634 -654 -1628
rect -735 -1659 -722 -1634
rect -691 -1659 -678 -1634
rect 1869 -1644 1889 -1640
rect 1900 -1644 1931 -1640
rect 1943 -1644 1971 -1640
rect 1981 -1644 2002 -1640
rect 2018 -1642 2048 -1638
rect 1869 -1647 1873 -1644
rect 1907 -1647 1911 -1644
rect 1951 -1647 1955 -1644
rect 1989 -1647 1993 -1644
rect 2035 -1645 2039 -1642
rect 1863 -1651 1864 -1647
rect 1868 -1651 1873 -1647
rect 1901 -1651 1902 -1647
rect 1906 -1651 1911 -1647
rect 1945 -1651 1946 -1647
rect 1950 -1651 1955 -1647
rect 1983 -1651 1984 -1647
rect 1988 -1651 1993 -1647
rect 2029 -1649 2030 -1645
rect 2034 -1649 2039 -1645
rect -796 -1670 -789 -1666
rect -785 -1678 -776 -1674
rect -769 -1681 -765 -1659
rect -761 -1670 -760 -1666
rect -725 -1668 -722 -1659
rect -681 -1668 -678 -1659
rect -725 -1673 -713 -1668
rect -681 -1673 -657 -1668
rect -650 -1669 -646 -1659
rect 1336 -1662 1340 -1654
rect 1364 -1662 1368 -1654
rect 1391 -1662 1395 -1654
rect 1430 -1662 1434 -1654
rect 1458 -1662 1462 -1654
rect 1485 -1662 1489 -1654
rect 1525 -1661 1529 -1653
rect 1553 -1661 1557 -1653
rect 1580 -1661 1584 -1653
rect 1616 -1661 1620 -1653
rect 1869 -1657 1873 -1651
rect 1907 -1657 1911 -1651
rect 1951 -1657 1955 -1651
rect 1989 -1657 1993 -1651
rect 2035 -1655 2039 -1649
rect -761 -1675 -753 -1673
rect -756 -1678 -753 -1675
rect -734 -1678 -733 -1674
rect -725 -1681 -722 -1673
rect -717 -1678 -709 -1673
rect -690 -1678 -689 -1674
rect -681 -1681 -678 -1673
rect -650 -1674 -637 -1669
rect -650 -1681 -646 -1674
rect -308 -1681 -280 -1678
rect -777 -1691 -765 -1681
rect -733 -1691 -722 -1681
rect -689 -1691 -678 -1681
rect -307 -1687 -304 -1681
rect -283 -1682 -280 -1681
rect -283 -1685 -212 -1682
rect -789 -1696 -785 -1691
rect -753 -1696 -749 -1691
rect -709 -1696 -705 -1691
rect -658 -1696 -654 -1691
rect -790 -1700 -646 -1696
rect -324 -1711 -321 -1708
rect -316 -1710 -306 -1707
rect -298 -1707 -295 -1699
rect -268 -1691 -265 -1685
rect -249 -1691 -246 -1685
rect -298 -1710 -277 -1707
rect -298 -1713 -295 -1710
rect -307 -1723 -304 -1719
rect -313 -1725 -289 -1723
rect -313 -1726 -295 -1725
rect -290 -1726 -289 -1725
rect -280 -1733 -277 -1710
rect -239 -1691 -219 -1688
rect -239 -1697 -236 -1691
rect -222 -1697 -219 -1691
rect -258 -1718 -255 -1715
rect -258 -1721 -240 -1718
rect -230 -1728 -227 -1721
rect -230 -1731 -213 -1728
rect -308 -1734 -289 -1733
rect -313 -1736 -289 -1734
rect -280 -1736 -237 -1733
rect -307 -1742 -304 -1736
rect -216 -1742 -213 -1731
rect -251 -1747 -226 -1744
rect -216 -1746 -203 -1742
rect -251 -1749 -248 -1747
rect -324 -1765 -321 -1762
rect -316 -1765 -306 -1762
rect -298 -1762 -295 -1754
rect -286 -1752 -248 -1749
rect -216 -1750 -213 -1746
rect -286 -1762 -283 -1752
rect -245 -1753 -213 -1750
rect -245 -1756 -242 -1753
rect -298 -1765 -283 -1762
rect -298 -1768 -295 -1765
rect -246 -1759 -240 -1756
rect -307 -1778 -304 -1774
rect -286 -1775 -281 -1772
rect -268 -1772 -265 -1768
rect -221 -1772 -218 -1768
rect -276 -1775 -212 -1772
rect -286 -1778 -283 -1775
rect -313 -1781 -283 -1778
rect -207 -1786 -203 -1746
rect 1877 -1715 1881 -1697
rect 1915 -1715 1919 -1697
rect 1959 -1715 1963 -1697
rect 1997 -1715 2001 -1697
rect 2043 -1713 2047 -1695
rect 1869 -1744 1873 -1735
rect 1907 -1744 1911 -1735
rect 1951 -1744 1955 -1735
rect 1989 -1744 1993 -1735
rect 2035 -1742 2039 -1733
rect 1869 -1748 1889 -1744
rect 1900 -1748 1931 -1744
rect 1943 -1748 1971 -1744
rect 1981 -1748 1998 -1744
rect 2018 -1746 2044 -1742
rect 1344 -1768 1348 -1762
rect 1372 -1768 1376 -1762
rect 1399 -1768 1403 -1762
rect 1438 -1768 1442 -1762
rect 1466 -1768 1470 -1762
rect 1493 -1768 1497 -1762
rect 1533 -1767 1537 -1761
rect 1561 -1767 1565 -1761
rect 1588 -1767 1592 -1761
rect 1624 -1767 1628 -1761
rect -787 -1790 -634 -1786
rect -781 -1796 -777 -1790
rect -743 -1796 -739 -1790
rect -699 -1796 -695 -1790
rect -654 -1796 -650 -1790
rect -731 -1821 -718 -1796
rect -687 -1821 -674 -1796
rect -792 -1832 -785 -1828
rect -781 -1840 -772 -1836
rect -765 -1843 -761 -1821
rect -757 -1832 -756 -1828
rect -721 -1830 -718 -1821
rect -677 -1830 -674 -1821
rect -721 -1835 -709 -1830
rect -677 -1835 -653 -1830
rect -646 -1831 -642 -1821
rect -757 -1837 -749 -1835
rect -752 -1840 -749 -1837
rect -730 -1840 -729 -1836
rect -721 -1843 -718 -1835
rect -713 -1840 -705 -1835
rect -686 -1840 -685 -1836
rect -677 -1843 -674 -1835
rect -646 -1836 -633 -1831
rect -646 -1843 -642 -1836
rect -773 -1853 -761 -1843
rect -729 -1853 -718 -1843
rect -685 -1853 -674 -1843
rect -785 -1858 -781 -1853
rect -749 -1858 -745 -1853
rect -705 -1858 -701 -1853
rect -654 -1858 -650 -1853
rect -786 -1862 -642 -1858
rect 4073 -1867 4226 -1863
rect 191 -1873 214 -1869
rect 195 -1875 214 -1873
rect 191 -1884 195 -1879
rect 210 -1884 214 -1875
rect 4079 -1873 4083 -1867
rect 4117 -1873 4121 -1867
rect 4161 -1873 4165 -1867
rect 4206 -1873 4210 -1867
rect 227 -1880 251 -1879
rect 227 -1884 243 -1880
rect 247 -1884 251 -1880
rect 227 -1886 251 -1884
rect 233 -1891 237 -1886
rect 202 -1912 206 -1904
rect 4129 -1898 4142 -1873
rect 4173 -1898 4186 -1873
rect 4068 -1909 4075 -1905
rect 202 -1916 214 -1912
rect 210 -1918 214 -1916
rect 241 -1918 245 -1911
rect 4079 -1917 4088 -1913
rect 185 -1923 203 -1919
rect 210 -1922 234 -1918
rect 241 -1922 251 -1918
rect 4095 -1920 4099 -1898
rect 4103 -1909 4104 -1905
rect 4139 -1907 4142 -1898
rect 4183 -1907 4186 -1898
rect 4139 -1912 4151 -1907
rect 4183 -1912 4207 -1907
rect 4214 -1908 4218 -1898
rect 4103 -1914 4111 -1912
rect 4108 -1917 4111 -1914
rect 4130 -1917 4131 -1913
rect 4139 -1920 4142 -1912
rect 4147 -1917 4155 -1912
rect 4174 -1917 4175 -1913
rect 4183 -1920 4186 -1912
rect 4214 -1913 4227 -1908
rect 4214 -1920 4218 -1913
rect 185 -1930 192 -1926
rect 210 -1933 214 -1922
rect 241 -1925 245 -1922
rect 4087 -1930 4099 -1920
rect 4131 -1930 4142 -1920
rect 4175 -1930 4186 -1920
rect 4075 -1935 4079 -1930
rect 4111 -1935 4115 -1930
rect 4155 -1935 4159 -1930
rect 4206 -1935 4210 -1930
rect 233 -1939 237 -1935
rect 4074 -1939 4218 -1935
rect 227 -1940 252 -1939
rect 227 -1944 247 -1940
rect 227 -1945 252 -1944
rect 191 -1957 195 -1953
rect 191 -1961 207 -1957
rect 3703 -1995 3731 -1992
rect 3704 -2001 3707 -1995
rect 3728 -1996 3731 -1995
rect 3728 -1999 3799 -1996
rect 3687 -2025 3690 -2022
rect 3695 -2024 3705 -2021
rect 3713 -2021 3716 -2013
rect 3743 -2005 3746 -1999
rect 3762 -2005 3765 -1999
rect 3713 -2024 3734 -2021
rect 3713 -2027 3716 -2024
rect -782 -2040 -629 -2036
rect 3704 -2037 3707 -2033
rect -281 -2040 -253 -2037
rect 3698 -2039 3722 -2037
rect 3698 -2040 3716 -2039
rect -776 -2046 -772 -2040
rect -738 -2046 -734 -2040
rect -694 -2046 -690 -2040
rect -649 -2046 -645 -2040
rect -280 -2046 -277 -2040
rect -256 -2041 -253 -2040
rect -256 -2044 -185 -2041
rect -726 -2071 -713 -2046
rect -682 -2071 -669 -2046
rect -297 -2070 -294 -2067
rect -289 -2069 -279 -2066
rect -271 -2066 -268 -2058
rect -241 -2050 -238 -2044
rect -222 -2050 -219 -2044
rect -271 -2069 -250 -2066
rect -787 -2082 -780 -2078
rect -776 -2090 -767 -2086
rect -760 -2093 -756 -2071
rect -752 -2082 -751 -2078
rect -716 -2080 -713 -2071
rect -672 -2080 -669 -2071
rect -716 -2085 -704 -2080
rect -672 -2085 -648 -2080
rect -641 -2081 -637 -2071
rect -271 -2072 -268 -2069
rect -752 -2087 -744 -2085
rect -747 -2090 -744 -2087
rect -725 -2090 -724 -2086
rect -716 -2093 -713 -2085
rect -708 -2090 -700 -2085
rect -681 -2090 -680 -2086
rect -672 -2093 -669 -2085
rect -641 -2086 -628 -2081
rect -280 -2082 -277 -2078
rect -286 -2084 -262 -2082
rect -286 -2085 -268 -2084
rect -641 -2093 -637 -2086
rect -768 -2103 -756 -2093
rect -724 -2103 -713 -2093
rect -680 -2103 -669 -2093
rect -263 -2085 -262 -2084
rect -253 -2092 -250 -2069
rect -212 -2050 -192 -2047
rect 3721 -2040 3722 -2039
rect 3731 -2047 3734 -2024
rect 3772 -2005 3792 -2002
rect 3772 -2011 3775 -2005
rect 3789 -2011 3792 -2005
rect 3753 -2032 3756 -2029
rect 3753 -2035 3771 -2032
rect 3781 -2042 3784 -2035
rect 3781 -2045 3798 -2042
rect 3703 -2048 3722 -2047
rect 3698 -2050 3722 -2048
rect 3731 -2050 3774 -2047
rect -212 -2056 -209 -2050
rect -195 -2056 -192 -2050
rect 3704 -2056 3707 -2050
rect 3795 -2056 3798 -2045
rect -231 -2077 -228 -2074
rect -231 -2080 -213 -2077
rect 3760 -2061 3785 -2058
rect 3795 -2060 3808 -2056
rect 3760 -2063 3763 -2061
rect 3687 -2079 3690 -2076
rect 3695 -2079 3705 -2076
rect 3713 -2076 3716 -2068
rect 3725 -2066 3763 -2063
rect 3795 -2064 3798 -2060
rect 3725 -2076 3728 -2066
rect 3766 -2067 3798 -2064
rect 3766 -2070 3769 -2067
rect 3713 -2079 3728 -2076
rect -203 -2087 -200 -2080
rect 3713 -2082 3716 -2079
rect -203 -2090 -186 -2087
rect -281 -2093 -262 -2092
rect -286 -2095 -262 -2093
rect -253 -2095 -210 -2092
rect -280 -2101 -277 -2095
rect -189 -2101 -186 -2090
rect 3765 -2073 3771 -2070
rect 3704 -2092 3707 -2088
rect 3725 -2089 3730 -2086
rect 3743 -2086 3746 -2082
rect 3790 -2086 3793 -2082
rect 3735 -2089 3799 -2086
rect 3725 -2092 3728 -2089
rect 3698 -2095 3728 -2092
rect 3804 -2100 3808 -2060
rect -780 -2108 -776 -2103
rect -744 -2108 -740 -2103
rect -700 -2108 -696 -2103
rect -649 -2108 -645 -2103
rect -781 -2112 -637 -2108
rect -224 -2106 -199 -2103
rect -189 -2105 -176 -2101
rect -224 -2108 -221 -2106
rect -297 -2124 -294 -2121
rect -289 -2124 -279 -2121
rect -271 -2121 -268 -2113
rect -259 -2111 -221 -2108
rect -189 -2109 -186 -2105
rect -259 -2121 -256 -2111
rect -218 -2112 -186 -2109
rect -218 -2115 -215 -2112
rect -271 -2124 -256 -2121
rect -271 -2127 -268 -2124
rect -219 -2118 -213 -2115
rect -280 -2137 -277 -2133
rect -259 -2134 -254 -2131
rect -241 -2131 -238 -2127
rect -194 -2131 -191 -2127
rect -249 -2134 -185 -2131
rect -259 -2137 -256 -2134
rect -286 -2140 -256 -2137
rect -180 -2145 -176 -2105
rect 199 -2165 222 -2161
rect 203 -2167 222 -2165
rect 199 -2176 203 -2171
rect 218 -2176 222 -2167
rect 235 -2172 259 -2171
rect 235 -2176 251 -2172
rect 255 -2176 259 -2172
rect 235 -2178 259 -2176
rect 241 -2183 245 -2178
rect -784 -2200 -631 -2196
rect -778 -2206 -774 -2200
rect -740 -2206 -736 -2200
rect -696 -2206 -692 -2200
rect -651 -2206 -647 -2200
rect 210 -2204 214 -2196
rect -728 -2231 -715 -2206
rect -684 -2231 -671 -2206
rect 210 -2208 222 -2204
rect 218 -2210 222 -2208
rect 249 -2210 253 -2203
rect 193 -2215 211 -2211
rect 218 -2214 242 -2210
rect 249 -2214 259 -2210
rect 193 -2222 200 -2218
rect 218 -2225 222 -2214
rect 249 -2217 253 -2214
rect -789 -2242 -782 -2238
rect -778 -2250 -769 -2246
rect -762 -2253 -758 -2231
rect -754 -2242 -753 -2238
rect -718 -2240 -715 -2231
rect -674 -2240 -671 -2231
rect -718 -2245 -706 -2240
rect -674 -2245 -650 -2240
rect -643 -2241 -639 -2231
rect -754 -2247 -746 -2245
rect -749 -2250 -746 -2247
rect -727 -2250 -726 -2246
rect -718 -2253 -715 -2245
rect -710 -2250 -702 -2245
rect -683 -2250 -682 -2246
rect -674 -2253 -671 -2245
rect -643 -2246 -630 -2241
rect 241 -2231 245 -2227
rect 235 -2232 260 -2231
rect 235 -2236 255 -2232
rect 235 -2237 260 -2236
rect -643 -2253 -639 -2246
rect 199 -2249 203 -2245
rect 199 -2253 215 -2249
rect -770 -2263 -758 -2253
rect -726 -2263 -715 -2253
rect -682 -2263 -671 -2253
rect -782 -2268 -778 -2263
rect -746 -2268 -742 -2263
rect -702 -2268 -698 -2263
rect -651 -2268 -647 -2263
rect -783 -2272 -639 -2268
rect -288 -2383 -260 -2380
rect -287 -2389 -284 -2383
rect -263 -2384 -260 -2383
rect -263 -2387 -192 -2384
rect -304 -2413 -301 -2410
rect -296 -2412 -286 -2409
rect -278 -2409 -275 -2401
rect -248 -2393 -245 -2387
rect -229 -2393 -226 -2387
rect -278 -2412 -257 -2409
rect -278 -2415 -275 -2412
rect -287 -2425 -284 -2421
rect -293 -2427 -269 -2425
rect -293 -2428 -275 -2427
rect -756 -2435 -603 -2431
rect -750 -2441 -746 -2435
rect -712 -2441 -708 -2435
rect -668 -2441 -664 -2435
rect -623 -2441 -619 -2435
rect -270 -2428 -269 -2427
rect -260 -2435 -257 -2412
rect -219 -2393 -199 -2390
rect -219 -2399 -216 -2393
rect -202 -2399 -199 -2393
rect -238 -2420 -235 -2417
rect -238 -2423 -220 -2420
rect 4058 -2420 4211 -2416
rect -210 -2430 -207 -2423
rect 3643 -2425 3671 -2422
rect -210 -2433 -193 -2430
rect -288 -2436 -269 -2435
rect -293 -2438 -269 -2436
rect -260 -2438 -217 -2435
rect -700 -2466 -687 -2441
rect -656 -2466 -643 -2441
rect -287 -2444 -284 -2438
rect -196 -2444 -193 -2433
rect 3644 -2431 3647 -2425
rect 3668 -2426 3671 -2425
rect 4064 -2426 4068 -2420
rect 4102 -2426 4106 -2420
rect 4146 -2426 4150 -2420
rect 4191 -2426 4195 -2420
rect 3668 -2429 3739 -2426
rect -231 -2449 -206 -2446
rect -196 -2448 -183 -2444
rect -231 -2451 -228 -2449
rect -761 -2477 -754 -2473
rect -750 -2485 -741 -2481
rect -734 -2488 -730 -2466
rect -726 -2477 -725 -2473
rect -690 -2475 -687 -2466
rect -646 -2475 -643 -2466
rect -690 -2480 -678 -2475
rect -646 -2480 -622 -2475
rect -615 -2476 -611 -2466
rect -304 -2467 -301 -2464
rect -296 -2467 -286 -2464
rect -278 -2464 -275 -2456
rect -266 -2454 -228 -2451
rect -196 -2452 -193 -2448
rect -266 -2464 -263 -2454
rect -225 -2455 -193 -2452
rect -225 -2458 -222 -2455
rect -278 -2467 -263 -2464
rect -278 -2470 -275 -2467
rect -226 -2461 -220 -2458
rect -726 -2482 -718 -2480
rect -721 -2485 -718 -2482
rect -699 -2485 -698 -2481
rect -690 -2488 -687 -2480
rect -682 -2485 -674 -2480
rect -655 -2485 -654 -2481
rect -646 -2488 -643 -2480
rect -615 -2481 -602 -2476
rect -287 -2480 -284 -2476
rect -266 -2477 -261 -2474
rect -248 -2474 -245 -2470
rect -201 -2474 -198 -2470
rect -256 -2477 -192 -2474
rect -266 -2480 -263 -2477
rect -615 -2488 -611 -2481
rect -293 -2483 -263 -2480
rect -187 -2488 -183 -2448
rect 3627 -2455 3630 -2452
rect 3635 -2454 3645 -2451
rect 3653 -2451 3656 -2443
rect 3683 -2435 3686 -2429
rect 3702 -2435 3705 -2429
rect 3653 -2454 3674 -2451
rect 3653 -2457 3656 -2454
rect 3644 -2467 3647 -2463
rect 3638 -2469 3662 -2467
rect 3638 -2470 3656 -2469
rect 3661 -2470 3662 -2469
rect 3671 -2477 3674 -2454
rect 3712 -2435 3732 -2432
rect 3712 -2441 3715 -2435
rect 3729 -2441 3732 -2435
rect 3693 -2462 3696 -2459
rect 3693 -2465 3711 -2462
rect 4114 -2451 4127 -2426
rect 4158 -2451 4171 -2426
rect 4053 -2462 4060 -2458
rect 3721 -2472 3724 -2465
rect 4064 -2470 4073 -2466
rect 3721 -2475 3738 -2472
rect 4080 -2473 4084 -2451
rect 4088 -2462 4089 -2458
rect 4124 -2460 4127 -2451
rect 4168 -2460 4171 -2451
rect 4124 -2465 4136 -2460
rect 4168 -2465 4192 -2460
rect 4199 -2461 4203 -2451
rect 4088 -2467 4096 -2465
rect 4093 -2470 4096 -2467
rect 4115 -2470 4116 -2466
rect 4124 -2473 4127 -2465
rect 4132 -2470 4140 -2465
rect 4159 -2470 4160 -2466
rect 4168 -2473 4171 -2465
rect 4199 -2466 4212 -2461
rect 4199 -2473 4203 -2466
rect 3643 -2478 3662 -2477
rect 3638 -2480 3662 -2478
rect 3671 -2480 3714 -2477
rect 3644 -2486 3647 -2480
rect 3735 -2486 3738 -2475
rect 4072 -2483 4084 -2473
rect 4116 -2483 4127 -2473
rect 4160 -2483 4171 -2473
rect -742 -2498 -730 -2488
rect -698 -2498 -687 -2488
rect -654 -2498 -643 -2488
rect 3700 -2491 3725 -2488
rect 3735 -2490 3748 -2486
rect 4060 -2488 4064 -2483
rect 4096 -2488 4100 -2483
rect 4140 -2488 4144 -2483
rect 4191 -2488 4195 -2483
rect 3700 -2493 3703 -2491
rect -754 -2503 -750 -2498
rect -718 -2503 -714 -2498
rect -674 -2503 -670 -2498
rect -623 -2503 -619 -2498
rect -755 -2507 -611 -2503
rect 3627 -2509 3630 -2506
rect 3635 -2509 3645 -2506
rect 3653 -2506 3656 -2498
rect 3665 -2496 3703 -2493
rect 3735 -2494 3738 -2490
rect 3665 -2506 3668 -2496
rect 3706 -2497 3738 -2494
rect 3706 -2500 3709 -2497
rect 3653 -2509 3668 -2506
rect 3653 -2512 3656 -2509
rect 3705 -2503 3711 -2500
rect 3644 -2522 3647 -2518
rect 3665 -2519 3670 -2516
rect 3683 -2516 3686 -2512
rect 3730 -2516 3733 -2512
rect 3675 -2519 3739 -2516
rect 3665 -2522 3668 -2519
rect 3638 -2525 3668 -2522
rect 187 -2531 210 -2527
rect 3744 -2530 3748 -2490
rect 4059 -2492 4203 -2488
rect 191 -2533 210 -2531
rect 187 -2542 191 -2537
rect 206 -2542 210 -2533
rect -747 -2560 -594 -2556
rect -741 -2566 -737 -2560
rect -703 -2566 -699 -2560
rect -659 -2566 -655 -2560
rect -614 -2566 -610 -2560
rect 223 -2538 247 -2537
rect 223 -2542 239 -2538
rect 243 -2542 247 -2538
rect 223 -2544 247 -2542
rect 229 -2549 233 -2544
rect -691 -2591 -678 -2566
rect -647 -2591 -634 -2566
rect 198 -2570 202 -2562
rect 198 -2574 210 -2570
rect 206 -2576 210 -2574
rect 237 -2576 241 -2569
rect 181 -2581 199 -2577
rect 206 -2580 230 -2576
rect 237 -2580 247 -2576
rect 181 -2588 188 -2584
rect 206 -2591 210 -2580
rect 237 -2583 241 -2580
rect -752 -2602 -745 -2598
rect -741 -2610 -732 -2606
rect -725 -2613 -721 -2591
rect -717 -2602 -716 -2598
rect -681 -2600 -678 -2591
rect -637 -2600 -634 -2591
rect -681 -2605 -669 -2600
rect -637 -2605 -613 -2600
rect -606 -2601 -602 -2591
rect -717 -2607 -709 -2605
rect -712 -2610 -709 -2607
rect -690 -2610 -689 -2606
rect -681 -2613 -678 -2605
rect -673 -2610 -665 -2605
rect -646 -2610 -645 -2606
rect -637 -2613 -634 -2605
rect -606 -2606 -593 -2601
rect -606 -2613 -602 -2606
rect -733 -2623 -721 -2613
rect -689 -2623 -678 -2613
rect -645 -2623 -634 -2613
rect 229 -2597 233 -2593
rect 223 -2598 248 -2597
rect 223 -2602 243 -2598
rect 223 -2603 248 -2602
rect 187 -2615 191 -2611
rect 187 -2619 203 -2615
rect -745 -2628 -741 -2623
rect -709 -2628 -705 -2623
rect -665 -2628 -661 -2623
rect -614 -2628 -610 -2623
rect -746 -2632 -602 -2628
rect 4071 -2712 4224 -2708
rect 4077 -2718 4081 -2712
rect 4115 -2718 4119 -2712
rect 4159 -2718 4163 -2712
rect 4204 -2718 4208 -2712
rect 4127 -2743 4140 -2718
rect 4171 -2743 4184 -2718
rect 4066 -2754 4073 -2750
rect 4077 -2762 4086 -2758
rect 4093 -2765 4097 -2743
rect 4101 -2754 4102 -2750
rect 4137 -2752 4140 -2743
rect 4181 -2752 4184 -2743
rect 4137 -2757 4149 -2752
rect 4181 -2757 4205 -2752
rect 4212 -2753 4216 -2743
rect 4101 -2759 4109 -2757
rect 4106 -2762 4109 -2759
rect 4128 -2762 4129 -2758
rect 4137 -2765 4140 -2757
rect 4145 -2762 4153 -2757
rect 4172 -2762 4173 -2758
rect 4181 -2765 4184 -2757
rect 4212 -2758 4225 -2753
rect 4212 -2765 4216 -2758
rect 4085 -2775 4097 -2765
rect 4129 -2775 4140 -2765
rect 4173 -2775 4184 -2765
rect 4073 -2780 4077 -2775
rect 4109 -2780 4113 -2775
rect 4153 -2780 4157 -2775
rect 4204 -2780 4208 -2775
rect 4072 -2784 4216 -2780
rect 3600 -2961 3628 -2958
rect 3601 -2967 3604 -2961
rect 3625 -2962 3628 -2961
rect 3625 -2965 3696 -2962
rect 3584 -2991 3587 -2988
rect 3592 -2990 3602 -2987
rect 3610 -2987 3613 -2979
rect 3640 -2971 3643 -2965
rect 3659 -2971 3662 -2965
rect 3610 -2990 3631 -2987
rect 3610 -2993 3613 -2990
rect 3601 -3003 3604 -2999
rect 3595 -3005 3619 -3003
rect 3595 -3006 3613 -3005
rect 3618 -3006 3619 -3005
rect 3628 -3013 3631 -2990
rect 3669 -2971 3689 -2968
rect 3669 -2977 3672 -2971
rect 3686 -2977 3689 -2971
rect 3650 -2998 3653 -2995
rect 3650 -3001 3668 -2998
rect 3678 -3008 3681 -3001
rect 3678 -3011 3695 -3008
rect 3600 -3014 3619 -3013
rect 3595 -3016 3619 -3014
rect 3628 -3016 3671 -3013
rect 3601 -3022 3604 -3016
rect 3692 -3022 3695 -3011
rect 3657 -3027 3682 -3024
rect 3692 -3026 3705 -3022
rect 3657 -3029 3660 -3027
rect 3584 -3045 3587 -3042
rect 3592 -3045 3602 -3042
rect 3610 -3042 3613 -3034
rect 3622 -3032 3660 -3029
rect 3692 -3030 3695 -3026
rect 3622 -3042 3625 -3032
rect 3663 -3033 3695 -3030
rect 3663 -3036 3666 -3033
rect 3610 -3045 3625 -3042
rect 3610 -3048 3613 -3045
rect 3662 -3039 3668 -3036
rect 3601 -3058 3604 -3054
rect 3622 -3055 3627 -3052
rect 3640 -3052 3643 -3048
rect 3687 -3052 3690 -3048
rect 3632 -3055 3696 -3052
rect 3622 -3058 3625 -3055
rect 3595 -3061 3625 -3058
rect 3701 -3066 3705 -3026
rect 4093 -3086 4246 -3082
rect 4099 -3092 4103 -3086
rect 4137 -3092 4141 -3086
rect 4181 -3092 4185 -3086
rect 4226 -3092 4230 -3086
rect 4149 -3117 4162 -3092
rect 4193 -3117 4206 -3092
rect 4088 -3128 4095 -3124
rect 4099 -3136 4108 -3132
rect 4115 -3139 4119 -3117
rect 4123 -3128 4124 -3124
rect 4159 -3126 4162 -3117
rect 4203 -3126 4206 -3117
rect 4159 -3131 4171 -3126
rect 4203 -3131 4227 -3126
rect 4234 -3127 4238 -3117
rect 4123 -3133 4131 -3131
rect 4128 -3136 4131 -3133
rect 4150 -3136 4151 -3132
rect 4159 -3139 4162 -3131
rect 4167 -3136 4175 -3131
rect 4194 -3136 4195 -3132
rect 4203 -3139 4206 -3131
rect 4234 -3132 4247 -3127
rect 4234 -3139 4238 -3132
rect 4107 -3149 4119 -3139
rect 4151 -3149 4162 -3139
rect 4195 -3149 4206 -3139
rect 4095 -3154 4099 -3149
rect 4131 -3154 4135 -3149
rect 4175 -3154 4179 -3149
rect 4226 -3154 4230 -3149
rect 4094 -3158 4238 -3154
<< m2contact >>
rect -832 -1013 -827 -1008
rect -802 -1005 -797 -1000
rect -803 -1015 -798 -1010
rect -775 -1013 -770 -1008
rect -731 -1013 -726 -1008
rect -838 -1182 -833 -1177
rect -808 -1174 -803 -1169
rect -809 -1184 -804 -1179
rect -781 -1182 -776 -1177
rect -737 -1182 -732 -1177
rect 3650 -1216 3655 -1211
rect 3650 -1270 3655 -1265
rect -838 -1362 -833 -1357
rect -808 -1354 -803 -1349
rect -312 -1353 -307 -1348
rect -809 -1364 -804 -1359
rect -781 -1362 -776 -1357
rect -737 -1362 -732 -1357
rect -312 -1407 -307 -1402
rect 4089 -1476 4094 -1471
rect 4119 -1468 4124 -1463
rect 4118 -1478 4123 -1473
rect 4146 -1476 4151 -1471
rect 4190 -1476 4195 -1471
rect -790 -1678 -785 -1673
rect -760 -1670 -755 -1665
rect -761 -1680 -756 -1675
rect -733 -1678 -728 -1673
rect -689 -1678 -684 -1673
rect -321 -1712 -316 -1707
rect -321 -1766 -316 -1761
rect -786 -1840 -781 -1835
rect -756 -1832 -751 -1827
rect -757 -1842 -752 -1837
rect -729 -1840 -724 -1835
rect -685 -1840 -680 -1835
rect 4074 -1917 4079 -1912
rect 4104 -1909 4109 -1904
rect 4103 -1919 4108 -1914
rect 4131 -1917 4136 -1912
rect 4175 -1917 4180 -1912
rect 3690 -2026 3695 -2021
rect -294 -2071 -289 -2066
rect -781 -2090 -776 -2085
rect -751 -2082 -746 -2077
rect -752 -2092 -747 -2087
rect -724 -2090 -719 -2085
rect -680 -2090 -675 -2085
rect 3690 -2080 3695 -2075
rect -294 -2125 -289 -2120
rect -783 -2250 -778 -2245
rect -753 -2242 -748 -2237
rect -754 -2252 -749 -2247
rect -726 -2250 -721 -2245
rect -682 -2250 -677 -2245
rect -301 -2414 -296 -2409
rect -755 -2485 -750 -2480
rect -725 -2477 -720 -2472
rect -301 -2468 -296 -2463
rect -726 -2487 -721 -2482
rect -698 -2485 -693 -2480
rect -654 -2485 -649 -2480
rect 3630 -2456 3635 -2451
rect 4059 -2470 4064 -2465
rect 4089 -2462 4094 -2457
rect 4088 -2472 4093 -2467
rect 4116 -2470 4121 -2465
rect 4160 -2470 4165 -2465
rect 3630 -2510 3635 -2505
rect -746 -2610 -741 -2605
rect -716 -2602 -711 -2597
rect -717 -2612 -712 -2607
rect -689 -2610 -684 -2605
rect -645 -2610 -640 -2605
rect 4072 -2762 4077 -2757
rect 4102 -2754 4107 -2749
rect 4101 -2764 4106 -2759
rect 4129 -2762 4134 -2757
rect 4173 -2762 4178 -2757
rect 3587 -2992 3592 -2987
rect 3587 -3046 3592 -3041
rect 4094 -3136 4099 -3131
rect 4124 -3128 4129 -3123
rect 4123 -3138 4128 -3133
rect 4151 -3136 4156 -3131
rect 4195 -3136 4200 -3131
<< pm12contact >>
rect 3706 -1233 3711 -1228
rect 3715 -1234 3720 -1229
rect -256 -1370 -251 -1365
rect -247 -1371 -242 -1366
rect 1399 -1499 1405 -1493
rect 1449 -1498 1455 -1492
rect 1499 -1498 1505 -1492
rect 1546 -1498 1552 -1492
rect -265 -1729 -260 -1724
rect -256 -1730 -251 -1725
rect 1869 -1712 1874 -1707
rect 1907 -1712 1912 -1707
rect 1951 -1712 1956 -1707
rect 1989 -1712 1994 -1707
rect 2035 -1710 2040 -1705
rect 1336 -1774 1341 -1769
rect 1364 -1774 1369 -1769
rect 1391 -1774 1396 -1769
rect 1430 -1774 1435 -1769
rect 1458 -1774 1463 -1769
rect 1485 -1774 1490 -1769
rect 1525 -1773 1530 -1768
rect 1553 -1773 1558 -1768
rect 1580 -1773 1585 -1768
rect 1616 -1773 1621 -1768
rect 3746 -2043 3751 -2038
rect 3755 -2044 3760 -2039
rect -238 -2088 -233 -2083
rect -229 -2089 -224 -2084
rect -245 -2431 -240 -2426
rect -236 -2432 -231 -2427
rect 3686 -2473 3691 -2468
rect 3695 -2474 3700 -2469
rect 3643 -3009 3648 -3004
rect 3652 -3010 3657 -3005
<< metal2 >>
rect -802 -955 -771 -952
rect -802 -1000 -798 -955
rect -775 -1008 -771 -955
rect -853 -1013 -832 -1009
rect -841 -1037 -835 -1013
rect -802 -1037 -798 -1015
rect -731 -1037 -726 -1013
rect -841 -1040 -722 -1037
rect -808 -1124 -777 -1121
rect -808 -1169 -804 -1124
rect -781 -1177 -777 -1124
rect -859 -1182 -838 -1178
rect -847 -1206 -841 -1182
rect -808 -1206 -804 -1184
rect -737 -1206 -732 -1182
rect -847 -1209 -728 -1206
rect 3651 -1222 3654 -1216
rect 3651 -1225 3688 -1222
rect 3685 -1228 3688 -1225
rect 3685 -1231 3706 -1228
rect 3715 -1244 3718 -1234
rect 3652 -1247 3718 -1244
rect 3652 -1265 3655 -1247
rect -808 -1304 -777 -1301
rect -808 -1349 -804 -1304
rect -781 -1357 -777 -1304
rect -859 -1362 -838 -1358
rect -847 -1386 -841 -1362
rect -311 -1359 -308 -1353
rect -311 -1362 -274 -1359
rect -808 -1386 -804 -1364
rect -737 -1386 -732 -1362
rect -277 -1365 -274 -1362
rect -277 -1368 -256 -1365
rect -247 -1381 -244 -1371
rect -310 -1384 -244 -1381
rect -847 -1389 -728 -1386
rect -310 -1402 -307 -1384
rect 4119 -1418 4150 -1415
rect 4119 -1463 4123 -1418
rect 4146 -1471 4150 -1418
rect 4068 -1476 4089 -1472
rect 1389 -1499 1399 -1493
rect 1439 -1498 1449 -1492
rect 1489 -1498 1499 -1492
rect 1536 -1498 1546 -1492
rect 4080 -1500 4086 -1476
rect 4119 -1500 4123 -1478
rect 4190 -1500 4195 -1476
rect 4080 -1503 4199 -1500
rect -760 -1620 -729 -1617
rect -760 -1665 -756 -1620
rect -733 -1673 -729 -1620
rect -811 -1678 -790 -1674
rect -799 -1702 -793 -1678
rect -760 -1702 -756 -1680
rect -689 -1702 -684 -1678
rect -799 -1705 -680 -1702
rect 1866 -1712 1869 -1707
rect 1904 -1712 1907 -1707
rect 1948 -1712 1951 -1707
rect 1986 -1712 1989 -1707
rect 2032 -1710 2035 -1705
rect -320 -1718 -317 -1712
rect -320 -1721 -283 -1718
rect -286 -1724 -283 -1721
rect -286 -1727 -265 -1724
rect -256 -1740 -253 -1730
rect -319 -1743 -253 -1740
rect -319 -1761 -316 -1743
rect 1332 -1774 1336 -1769
rect 1360 -1774 1364 -1769
rect 1387 -1774 1391 -1769
rect 1426 -1774 1430 -1769
rect 1454 -1774 1458 -1769
rect 1481 -1774 1485 -1769
rect 1521 -1773 1525 -1768
rect 1549 -1773 1553 -1768
rect 1576 -1773 1580 -1768
rect 1612 -1773 1616 -1768
rect -756 -1782 -725 -1779
rect -756 -1827 -752 -1782
rect -729 -1835 -725 -1782
rect -807 -1840 -786 -1836
rect -795 -1864 -789 -1840
rect -756 -1864 -752 -1842
rect -685 -1864 -680 -1840
rect 4104 -1859 4135 -1856
rect -795 -1867 -676 -1864
rect 4104 -1904 4108 -1859
rect 4131 -1912 4135 -1859
rect 4053 -1917 4074 -1913
rect 4065 -1941 4071 -1917
rect 4104 -1941 4108 -1919
rect 4175 -1941 4180 -1917
rect 4065 -1944 4184 -1941
rect -751 -2032 -720 -2029
rect -751 -2077 -747 -2032
rect -724 -2085 -720 -2032
rect 3691 -2032 3694 -2026
rect 3691 -2035 3728 -2032
rect 3725 -2038 3728 -2035
rect 3725 -2041 3746 -2038
rect 3755 -2054 3758 -2044
rect 3692 -2057 3758 -2054
rect -293 -2077 -290 -2071
rect 3692 -2075 3695 -2057
rect -293 -2080 -256 -2077
rect -259 -2083 -256 -2080
rect -802 -2090 -781 -2086
rect -790 -2114 -784 -2090
rect -751 -2114 -747 -2092
rect -680 -2114 -675 -2090
rect -259 -2086 -238 -2083
rect -229 -2099 -226 -2089
rect -292 -2102 -226 -2099
rect -790 -2117 -671 -2114
rect -292 -2120 -289 -2102
rect -753 -2192 -722 -2189
rect -753 -2237 -749 -2192
rect -726 -2245 -722 -2192
rect -804 -2250 -783 -2246
rect -792 -2274 -786 -2250
rect -753 -2274 -749 -2252
rect -682 -2274 -677 -2250
rect -792 -2277 -673 -2274
rect 4089 -2412 4120 -2409
rect -300 -2420 -297 -2414
rect -300 -2423 -263 -2420
rect -725 -2427 -694 -2424
rect -266 -2426 -263 -2423
rect -725 -2472 -721 -2427
rect -698 -2480 -694 -2427
rect -266 -2429 -245 -2426
rect -236 -2442 -233 -2432
rect -299 -2445 -233 -2442
rect -299 -2463 -296 -2445
rect 3631 -2462 3634 -2456
rect 4089 -2457 4093 -2412
rect 3631 -2465 3668 -2462
rect 4116 -2465 4120 -2412
rect 3665 -2468 3668 -2465
rect 3665 -2471 3686 -2468
rect 4038 -2470 4059 -2466
rect -776 -2485 -755 -2481
rect -764 -2509 -758 -2485
rect 3695 -2484 3698 -2474
rect -725 -2509 -721 -2487
rect -654 -2509 -649 -2485
rect 3632 -2487 3698 -2484
rect 3632 -2505 3635 -2487
rect 4050 -2494 4056 -2470
rect 4089 -2494 4093 -2472
rect 4160 -2494 4165 -2470
rect 4050 -2497 4169 -2494
rect -764 -2512 -645 -2509
rect -716 -2552 -685 -2549
rect -716 -2597 -712 -2552
rect -689 -2605 -685 -2552
rect -767 -2610 -746 -2606
rect -755 -2634 -749 -2610
rect -716 -2634 -712 -2612
rect -645 -2634 -640 -2610
rect -755 -2637 -636 -2634
rect 4102 -2704 4133 -2701
rect 4102 -2749 4106 -2704
rect 4129 -2757 4133 -2704
rect 4051 -2762 4072 -2758
rect 4063 -2786 4069 -2762
rect 4102 -2786 4106 -2764
rect 4173 -2786 4178 -2762
rect 4063 -2789 4182 -2786
rect 3588 -2998 3591 -2992
rect 3588 -3001 3625 -2998
rect 3622 -3004 3625 -3001
rect 3622 -3007 3643 -3004
rect 3652 -3020 3655 -3010
rect 3589 -3023 3655 -3020
rect 3589 -3041 3592 -3023
rect 4124 -3078 4155 -3075
rect 4124 -3123 4128 -3078
rect 4151 -3131 4155 -3078
rect 4073 -3136 4094 -3132
rect 4085 -3160 4091 -3136
rect 4124 -3160 4128 -3138
rect 4195 -3160 4200 -3136
rect 4085 -3163 4204 -3160
<< m123contact >>
rect 3658 -1185 3663 -1180
rect 3658 -1238 3663 -1233
rect 3676 -1234 3681 -1229
rect 3690 -1279 3695 -1274
rect -304 -1322 -299 -1317
rect -304 -1375 -299 -1370
rect -286 -1371 -281 -1366
rect -272 -1416 -267 -1411
rect -313 -1681 -308 -1676
rect -313 -1734 -308 -1729
rect -295 -1730 -290 -1725
rect -281 -1775 -276 -1770
rect 3698 -1995 3703 -1990
rect -286 -2040 -281 -2035
rect 3698 -2048 3703 -2043
rect 3716 -2044 3721 -2039
rect -286 -2093 -281 -2088
rect -268 -2089 -263 -2084
rect 3730 -2089 3735 -2084
rect -254 -2134 -249 -2129
rect -293 -2383 -288 -2378
rect 3638 -2425 3643 -2420
rect -293 -2436 -288 -2431
rect -275 -2432 -270 -2427
rect -261 -2477 -256 -2472
rect 3638 -2478 3643 -2473
rect 3656 -2474 3661 -2469
rect 3670 -2519 3675 -2514
rect 3595 -2961 3600 -2956
rect 3595 -3014 3600 -3009
rect 3613 -3010 3618 -3005
rect 3627 -3055 3632 -3050
<< metal3 >>
rect 3658 -1233 3661 -1185
rect 3681 -1234 3693 -1231
rect 3690 -1274 3693 -1234
rect -304 -1370 -301 -1322
rect -281 -1371 -269 -1368
rect -272 -1411 -269 -1371
rect -313 -1729 -310 -1681
rect -290 -1730 -278 -1727
rect -281 -1770 -278 -1730
rect -286 -2088 -283 -2040
rect 3698 -2043 3701 -1995
rect 3721 -2044 3733 -2041
rect 3730 -2084 3733 -2044
rect -263 -2089 -251 -2086
rect -254 -2129 -251 -2089
rect -293 -2431 -290 -2383
rect -270 -2432 -258 -2429
rect -261 -2472 -258 -2432
rect 3638 -2473 3641 -2425
rect 3661 -2474 3673 -2471
rect 3670 -2514 3673 -2474
rect 3595 -3009 3598 -2961
rect 3618 -3010 3630 -3007
rect 3627 -3050 3630 -3010
<< labels >>
rlabel metal1 1336 -1658 1340 -1654 1 pdr1
rlabel metal2 1332 -1774 1336 -1769 2 prop_1
rlabel metal1 1344 -1768 1348 -1763 1 prop1_car0
rlabel metal1 1364 -1659 1368 -1654 1 prop1_car0
rlabel metal2 1360 -1774 1364 -1769 1 carry_0
rlabel metal1 1372 -1768 1376 -1763 1 clock_car0
rlabel metal1 1391 -1659 1395 -1654 1 clock_car0
rlabel metal2 1387 -1774 1391 -1769 1 clock_in
rlabel metal1 1399 -1768 1403 -1763 1 gnd!
rlabel metal1 1430 -1659 1434 -1654 1 pdr2
rlabel metal2 1426 -1774 1430 -1769 1 prop_2
rlabel metal1 1438 -1768 1442 -1763 1 pdr1
rlabel metal1 1458 -1659 1462 -1654 1 pdr1
rlabel metal2 1454 -1774 1458 -1769 1 gen_1
rlabel metal1 1466 -1768 1470 -1763 1 clock_car0
rlabel metal1 1485 -1659 1489 -1654 1 pdr3
rlabel metal2 1481 -1774 1485 -1769 1 prop_3
rlabel metal1 1493 -1768 1497 -1763 1 pdr2
rlabel metal1 1525 -1658 1529 -1653 1 pdr2
rlabel metal2 1521 -1773 1525 -1768 1 gen_2
rlabel metal1 1533 -1767 1537 -1762 1 clock_car0
rlabel metal1 1553 -1658 1557 -1653 1 pdr4
rlabel metal2 1549 -1773 1553 -1768 1 prop_4
rlabel metal1 1561 -1767 1565 -1762 1 pdr3
rlabel metal1 1580 -1658 1584 -1653 1 pdr3
rlabel metal2 1576 -1773 1580 -1768 1 gen_3
rlabel metal1 1588 -1767 1592 -1762 1 clock_car0
rlabel metal1 1616 -1658 1620 -1653 1 pdr4
rlabel metal2 1612 -1773 1616 -1768 1 gen_4
rlabel metal1 1624 -1767 1628 -1762 7 clock_car0
rlabel metal1 1400 -1411 1404 -1406 5 vdd!
rlabel metal1 1450 -1410 1454 -1405 5 vdd!
rlabel metal1 1500 -1410 1504 -1405 5 vdd!
rlabel metal1 1547 -1410 1551 -1405 5 vdd!
rlabel metal2 1389 -1499 1395 -1493 2 clock_in
rlabel metal2 1439 -1498 1445 -1492 1 clock_in
rlabel metal2 1489 -1498 1495 -1492 1 clock_in
rlabel metal2 1536 -1498 1541 -1492 1 clock_in
rlabel metal1 1408 -1490 1412 -1485 1 pdr1
rlabel metal1 1458 -1489 1462 -1485 1 pdr2
rlabel metal1 1508 -1489 1512 -1485 1 pdr3
rlabel metal1 1555 -1489 1559 -1485 1 pdr4
rlabel metal1 1994 -1748 1998 -1744 1 gnd!
rlabel metal1 1990 -1644 1995 -1640 5 vdd!
rlabel metal2 1866 -1712 1869 -1707 1 pdr1
rlabel metal2 1904 -1712 1907 -1707 1 pdr2
rlabel metal2 1948 -1712 1951 -1707 1 pdr3
rlabel metal2 1986 -1712 1989 -1707 1 pdr4
rlabel metal1 1877 -1712 1881 -1707 1 c1
rlabel metal1 1915 -1712 1919 -1707 1 c2
rlabel metal1 1959 -1712 1963 -1707 1 c3
rlabel metal1 1997 -1712 2001 -1707 1 c4
rlabel metal1 2040 -1746 2044 -1742 1 gnd!
rlabel metal1 2036 -1642 2041 -1638 5 vdd!
rlabel metal2 2032 -1710 2035 -1705 1 clk_org
rlabel metal1 2043 -1710 2047 -1705 1 clock_in
rlabel metal1 1869 -1644 1873 -1640 5 vdd!
rlabel metal1 1907 -1644 1911 -1640 5 vdd!
rlabel metal1 1951 -1644 1955 -1640 5 vdd!
rlabel metal1 1955 -1748 1959 -1744 1 gnd!
rlabel metal1 1918 -1748 1922 -1744 1 gnd!
rlabel metal1 1878 -1748 1882 -1744 1 gnd!
rlabel metal1 199 -1522 199 -1522 5 vdd
rlabel metal1 200 -1609 200 -1609 1 gnd
rlabel metal1 232 -1591 232 -1591 1 gnd
rlabel metal1 229 -1534 229 -1534 5 vdd
rlabel metal1 201 -1872 201 -1872 5 vdd
rlabel metal1 202 -1959 202 -1959 1 gnd
rlabel metal1 234 -1941 234 -1941 1 gnd
rlabel metal1 231 -1884 231 -1884 5 vdd
rlabel metal1 209 -2164 209 -2164 5 vdd
rlabel metal1 210 -2251 210 -2251 1 gnd
rlabel metal1 242 -2233 242 -2233 1 gnd
rlabel metal1 239 -2176 239 -2176 5 vdd
rlabel metal1 197 -2530 197 -2530 5 vdd
rlabel metal1 198 -2617 198 -2617 1 gnd
rlabel metal1 230 -2599 230 -2599 1 gnd
rlabel metal1 227 -2542 227 -2542 5 vdd
rlabel metal1 184 -1571 184 -1571 3 q_a1
rlabel metal1 186 -1578 186 -1578 3 q_b1
rlabel metal1 248 -1571 248 -1571 1 gen_1
rlabel metal1 187 -1922 187 -1922 1 q_a2
rlabel metal1 187 -1929 187 -1929 1 q_b2
rlabel metal1 250 -1920 250 -1920 1 gen_2
rlabel metal1 194 -2214 194 -2214 1 q_b3
rlabel metal1 196 -2221 196 -2221 1 q_a3
rlabel metal1 257 -2212 257 -2212 1 gen_3
rlabel metal1 182 -2579 182 -2579 3 q_a4
rlabel metal1 182 -2585 182 -2585 3 q_b4
rlabel metal1 245 -2578 245 -2578 1 gen_4
rlabel metal1 -286 -1422 -282 -1419 1 gnd
rlabel metal1 -236 -1416 -233 -1414 1 gnd
rlabel metal1 -288 -1366 -287 -1364 1 gnd
rlabel metal1 -292 -1322 -289 -1320 5 vdd
rlabel metal1 -291 -1376 -288 -1374 1 vdd
rlabel metal1 -295 -1781 -291 -1778 1 gnd
rlabel metal1 -245 -1775 -242 -1773 1 gnd
rlabel metal1 -297 -1725 -296 -1723 1 gnd
rlabel metal1 -301 -1681 -298 -1679 5 vdd
rlabel metal1 -300 -1735 -297 -1733 1 vdd
rlabel metal1 -268 -2140 -264 -2137 1 gnd
rlabel metal1 -218 -2134 -215 -2132 1 gnd
rlabel metal1 -270 -2084 -269 -2082 1 gnd
rlabel metal1 -274 -2040 -271 -2038 5 vdd
rlabel metal1 -273 -2094 -270 -2092 1 vdd
rlabel metal1 -275 -2483 -271 -2480 1 gnd
rlabel metal1 -225 -2477 -222 -2475 1 gnd
rlabel metal1 -277 -2427 -276 -2425 1 gnd
rlabel metal1 -281 -2383 -278 -2381 5 vdd
rlabel metal1 -280 -2437 -277 -2435 1 vdd
rlabel metal1 3676 -1285 3680 -1282 1 gnd
rlabel metal1 3726 -1279 3729 -1277 1 gnd
rlabel metal1 3674 -1229 3675 -1227 1 gnd
rlabel metal1 3670 -1185 3673 -1183 5 vdd
rlabel metal1 3671 -1239 3674 -1237 1 vdd
rlabel metal1 3716 -2095 3720 -2092 1 gnd
rlabel metal1 3766 -2089 3769 -2087 1 gnd
rlabel metal1 3714 -2039 3715 -2037 1 gnd
rlabel metal1 3710 -1995 3713 -1993 5 vdd
rlabel metal1 3711 -2049 3714 -2047 1 vdd
rlabel metal1 3656 -2525 3660 -2522 1 gnd
rlabel metal1 3706 -2519 3709 -2517 1 gnd
rlabel metal1 3654 -2469 3655 -2467 1 gnd
rlabel metal1 3650 -2425 3653 -2423 5 vdd
rlabel metal1 3651 -2479 3654 -2477 1 vdd
rlabel metal1 -314 -1350 -314 -1350 1 q_a1
rlabel metal1 -314 -1404 -314 -1404 1 q_b1
rlabel metal1 -198 -1385 -198 -1385 1 prop_1
rlabel metal1 -323 -1709 -323 -1709 3 q_a2
rlabel metal1 -323 -1764 -323 -1764 3 q_b2
rlabel metal1 -205 -1743 -205 -1743 1 prop_2
rlabel metal1 -295 -2068 -295 -2068 1 q_a3
rlabel metal1 -295 -2122 -295 -2122 1 q_b3
rlabel metal1 -178 -2103 -178 -2103 1 prop_3
rlabel metal1 -303 -2412 -303 -2412 1 q_a4
rlabel metal1 -303 -2465 -303 -2465 1 q_b4
rlabel metal1 -184 -2446 -184 -2446 1 prop_4
rlabel metal1 3648 -1213 3648 -1213 1 carry_0
rlabel metal1 3648 -1267 3648 -1267 1 prop_1
rlabel metal1 3767 -1248 3767 -1248 1 s1
rlabel metal1 3689 -2024 3689 -2024 1 c1
rlabel metal1 3688 -2078 3688 -2078 1 prop_2
rlabel metal1 3807 -2059 3807 -2059 7 s2
rlabel metal1 3628 -2453 3628 -2453 1 c2
rlabel metal1 3628 -2508 3628 -2508 1 prop_3
rlabel metal1 3747 -2488 3747 -2488 1 s3
rlabel metal1 3613 -3061 3617 -3058 1 gnd
rlabel metal1 3663 -3055 3666 -3053 1 gnd
rlabel metal1 3611 -3005 3612 -3003 1 gnd
rlabel metal1 3607 -2961 3610 -2959 5 vdd
rlabel metal1 3608 -3015 3611 -3013 1 vdd
rlabel metal1 3703 -3024 3703 -3024 1 s4
rlabel metal1 3585 -3043 3585 -3043 1 prop_4
rlabel metal1 3585 -2990 3585 -2990 1 c3
rlabel metal1 -829 -1202 -826 -1201 1 gnd
rlabel metal1 -823 -1130 -821 -1129 5 vdd
rlabel metal2 -842 -1181 -842 -1181 1 clk_org
rlabel metal1 -829 -1382 -826 -1381 1 gnd
rlabel metal1 -823 -1310 -821 -1309 5 vdd
rlabel metal2 -842 -1361 -842 -1361 1 clk_org
rlabel metal1 -823 -1033 -820 -1032 1 gnd
rlabel metal1 -817 -961 -815 -960 5 vdd
rlabel metal2 -836 -1012 -836 -1012 1 clk_org
rlabel metal1 -781 -1698 -778 -1697 1 gnd
rlabel metal1 -775 -1626 -773 -1625 5 vdd
rlabel metal2 -794 -1677 -794 -1677 1 clk_org
rlabel metal1 -777 -1860 -774 -1859 1 gnd
rlabel metal1 -771 -1788 -769 -1787 5 vdd
rlabel metal2 -790 -1839 -790 -1839 1 clk_org
rlabel metal1 -772 -2110 -769 -2109 1 gnd
rlabel metal1 -766 -2038 -764 -2037 5 vdd
rlabel metal2 -785 -2089 -785 -2089 1 clk_org
rlabel metal1 -774 -2270 -771 -2269 1 gnd
rlabel metal1 -768 -2198 -766 -2197 5 vdd
rlabel metal2 -787 -2249 -787 -2249 1 clk_org
rlabel metal1 -746 -2505 -743 -2504 1 gnd
rlabel metal1 -740 -2433 -738 -2432 5 vdd
rlabel metal2 -759 -2484 -759 -2484 1 clk_org
rlabel metal1 -737 -2630 -734 -2629 1 gnd
rlabel metal1 -731 -2558 -729 -2557 5 vdd
rlabel metal2 -750 -2609 -750 -2609 1 clk_org
rlabel metal1 -837 -1003 -837 -1003 1 cin
rlabel metal1 -680 -1007 -680 -1007 1 carry_0
rlabel metal1 -842 -1172 -842 -1172 1 a1
rlabel metal1 -687 -1175 -687 -1175 1 q_a1
rlabel metal1 -842 -1352 -842 -1352 1 b1
rlabel metal1 -687 -1355 -687 -1355 1 q_b1
rlabel metal1 -794 -1668 -794 -1668 1 a2
rlabel metal1 -639 -1672 -639 -1672 1 q_a2
rlabel metal1 -789 -1830 -789 -1830 1 b2
rlabel metal1 -636 -1834 -636 -1834 1 q_b2
rlabel metal1 -785 -2080 -785 -2080 1 a3
rlabel metal1 -631 -2084 -631 -2084 1 q_a3
rlabel metal1 -786 -2240 -786 -2240 1 b3
rlabel metal1 -631 -2243 -631 -2243 1 q_b3
rlabel metal1 -759 -2474 -759 -2474 1 a4
rlabel metal1 -604 -2479 -604 -2479 1 q_a4
rlabel metal1 -750 -2600 -750 -2600 1 b4
rlabel metal1 -595 -2603 -595 -2603 1 q_b4
rlabel metal1 4098 -1496 4101 -1495 1 gnd
rlabel metal1 4104 -1424 4106 -1423 5 vdd
rlabel metal2 4085 -1475 4085 -1475 1 clk_org
rlabel metal1 4083 -1937 4086 -1936 1 gnd
rlabel metal1 4089 -1865 4091 -1864 5 vdd
rlabel metal2 4070 -1916 4070 -1916 1 clk_org
rlabel metal1 4068 -2490 4071 -2489 1 gnd
rlabel metal1 4074 -2418 4076 -2417 5 vdd
rlabel metal2 4055 -2469 4055 -2469 1 clk_org
rlabel metal1 4081 -2782 4084 -2781 1 gnd
rlabel metal1 4087 -2710 4089 -2709 5 vdd
rlabel metal2 4068 -2761 4068 -2761 1 clk_org
rlabel metal1 4085 -1466 4085 -1466 1 s1
rlabel metal1 4240 -1469 4240 -1469 7 q_s1
rlabel metal1 4071 -1907 4071 -1907 1 s2
rlabel metal1 4224 -1911 4224 -1911 1 q_s2
rlabel metal1 4055 -2460 4055 -2460 1 s3
rlabel metal1 4210 -2463 4210 -2463 1 q_s3
rlabel metal1 4068 -2752 4068 -2752 1 s4
rlabel metal1 4222 -2756 4222 -2756 1 q_s4
rlabel metal1 4103 -3156 4106 -3155 1 gnd
rlabel metal1 4109 -3084 4111 -3083 5 vdd
rlabel metal2 4090 -3135 4090 -3135 1 clk_org
rlabel metal1 4090 -3126 4090 -3126 1 c4
rlabel metal1 4245 -3129 4245 -3129 7 q_c4
<< end >>
