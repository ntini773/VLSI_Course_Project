magic
tech scmos
timestamp 1731964016
<< nwell >>
rect 6 35 39 82
rect 72 39 104 77
<< ntransistor >>
rect 22 17 24 27
rect 86 8 88 18
rect 77 -44 79 -34
<< ptransistor >>
rect 22 47 24 67
rect 86 50 88 70
<< ndiffusion >>
rect 21 17 22 27
rect 24 17 25 27
rect 85 8 86 18
rect 88 8 89 18
rect 76 -44 77 -34
rect 79 -44 80 -34
<< pdiffusion >>
rect 21 47 22 67
rect 24 47 25 67
rect 85 50 86 70
rect 88 50 89 70
<< ndcontact >>
rect 17 17 21 27
rect 25 17 29 27
rect 81 8 85 18
rect 89 8 93 18
rect 72 -44 76 -34
rect 80 -44 84 -34
<< pdcontact >>
rect 17 47 21 67
rect 25 47 29 67
rect 81 50 85 70
rect 89 50 93 70
<< polysilicon >>
rect 22 67 24 76
rect 86 70 88 80
rect 22 27 24 47
rect 86 35 88 50
rect 86 18 88 23
rect 22 14 24 17
rect 86 3 88 8
rect 77 -34 79 -13
rect 77 -51 79 -44
<< polycontact >>
rect 82 80 88 87
rect 18 30 22 34
rect 82 -4 88 3
rect 75 -13 79 -9
<< metal1 >>
rect -17 92 57 97
rect -17 -35 -11 92
rect 6 82 39 89
rect 53 87 57 92
rect 17 67 21 82
rect 53 80 82 87
rect -5 34 2 37
rect -5 30 18 34
rect 25 33 29 47
rect 53 34 60 80
rect 52 33 60 34
rect -5 -17 0 30
rect 25 29 60 33
rect 81 31 85 50
rect 25 27 29 29
rect 64 25 85 31
rect 81 18 85 25
rect 17 12 21 17
rect 6 5 42 12
rect 89 32 93 50
rect 89 26 124 32
rect 89 18 93 26
rect 56 -4 82 3
rect 56 -17 63 -4
rect -5 -23 63 -17
rect 67 -13 75 -9
rect 67 -27 70 -13
rect 118 -17 124 26
rect 64 -31 70 -27
rect 80 -23 124 -17
rect 64 -35 67 -31
rect 80 -34 84 -23
rect -17 -39 67 -35
rect 72 -57 76 -44
rect 60 -62 96 -57
<< labels >>
rlabel metal1 44 31 44 31 1 invo
rlabel metal1 8 32 8 32 1 invi
rlabel metal1 25 86 25 86 5 vdd
rlabel metal1 26 8 26 8 1 gnd
<< end >>
