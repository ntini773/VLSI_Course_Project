magic
tech scmos
timestamp 1733166931
<< nwell >>
rect -282 -111 -250 -74
rect -244 -111 -218 -74
rect -200 -111 -174 -74
rect -155 -111 -129 -74
<< ntransistor >>
rect -275 -137 -273 -127
rect -239 -137 -237 -127
rect -231 -137 -229 -127
rect -195 -137 -193 -127
rect -187 -137 -185 -127
rect -144 -137 -142 -127
<< ptransistor >>
rect -271 -105 -269 -80
rect -263 -105 -261 -80
rect -233 -105 -231 -80
rect -189 -105 -187 -80
rect -144 -105 -142 -80
<< ndiffusion >>
rect -276 -137 -275 -127
rect -273 -137 -272 -127
rect -240 -137 -239 -127
rect -237 -137 -236 -127
rect -232 -137 -231 -127
rect -229 -137 -228 -127
rect -196 -137 -195 -127
rect -193 -137 -192 -127
rect -188 -137 -187 -127
rect -185 -137 -184 -127
rect -145 -137 -144 -127
rect -142 -137 -141 -127
<< pdiffusion >>
rect -272 -105 -271 -80
rect -269 -105 -268 -80
rect -264 -105 -263 -80
rect -261 -105 -260 -80
rect -234 -105 -233 -80
rect -231 -105 -230 -80
rect -190 -105 -189 -80
rect -187 -105 -186 -80
rect -145 -105 -144 -80
rect -142 -105 -141 -80
<< ndcontact >>
rect -280 -137 -276 -127
rect -272 -137 -268 -127
rect -244 -137 -240 -127
rect -236 -137 -232 -127
rect -228 -137 -224 -127
rect -200 -137 -196 -127
rect -192 -137 -188 -127
rect -184 -137 -180 -127
rect -149 -137 -145 -127
rect -141 -137 -137 -127
<< pdcontact >>
rect -276 -105 -272 -80
rect -268 -105 -264 -80
rect -260 -105 -256 -80
rect -238 -105 -234 -80
rect -230 -105 -226 -80
rect -194 -105 -190 -80
rect -186 -105 -182 -80
rect -149 -105 -145 -80
rect -141 -105 -137 -80
<< polysilicon >>
rect -271 -80 -269 -77
rect -263 -80 -261 -77
rect -233 -80 -231 -77
rect -189 -80 -187 -77
rect -144 -80 -142 -77
rect -271 -112 -269 -105
rect -276 -116 -269 -112
rect -275 -127 -273 -116
rect -263 -124 -261 -105
rect -233 -113 -231 -105
rect -189 -113 -187 -105
rect -239 -115 -231 -113
rect -195 -115 -187 -113
rect -239 -127 -237 -115
rect -231 -127 -229 -118
rect -195 -127 -193 -115
rect -187 -127 -185 -118
rect -144 -127 -142 -105
rect -275 -140 -273 -137
rect -239 -140 -237 -137
rect -231 -140 -229 -137
rect -195 -140 -193 -137
rect -187 -140 -185 -137
rect -144 -140 -142 -137
<< polycontact >>
rect -280 -116 -276 -112
rect -267 -124 -263 -120
rect -256 -116 -252 -112
rect -244 -124 -239 -119
rect -229 -124 -225 -120
rect -200 -124 -195 -119
rect -148 -119 -144 -114
rect -185 -124 -181 -120
<< metal1 >>
rect -282 -74 -129 -70
rect -276 -80 -272 -74
rect -238 -80 -234 -74
rect -194 -80 -190 -74
rect -149 -80 -145 -74
rect -226 -105 -213 -80
rect -182 -105 -169 -80
rect -287 -116 -280 -112
rect -276 -124 -267 -120
rect -260 -127 -256 -105
rect -252 -116 -251 -112
rect -216 -114 -213 -105
rect -172 -114 -169 -105
rect -216 -119 -204 -114
rect -172 -119 -148 -114
rect -141 -115 -137 -105
rect -252 -121 -244 -119
rect -247 -124 -244 -121
rect -225 -124 -224 -120
rect -216 -127 -213 -119
rect -208 -124 -200 -119
rect -181 -124 -180 -120
rect -172 -127 -169 -119
rect -141 -120 -128 -115
rect -141 -127 -137 -120
rect -268 -137 -256 -127
rect -224 -137 -213 -127
rect -180 -137 -169 -127
rect -280 -142 -276 -137
rect -244 -142 -240 -137
rect -200 -142 -196 -137
rect -149 -142 -145 -137
rect -281 -146 -137 -142
<< m2contact >>
rect -281 -124 -276 -119
rect -251 -116 -246 -111
rect -252 -126 -247 -121
rect -224 -124 -219 -119
rect -180 -124 -175 -119
<< metal2 >>
rect -251 -66 -220 -63
rect -251 -111 -247 -66
rect -224 -119 -220 -66
rect -302 -124 -281 -120
rect -290 -148 -284 -124
rect -251 -148 -247 -126
rect -180 -148 -175 -124
rect -290 -151 -171 -148
<< labels >>
rlabel metal1 -272 -144 -269 -143 1 gnd
rlabel metal1 -266 -72 -264 -71 5 vdd
rlabel metal2 -285 -123 -285 -123 1 clk_org
rlabel metal1 -286 -114 -286 -114 1 a1
rlabel metal1 -129 -117 -129 -117 7 q_a1
<< end >>
