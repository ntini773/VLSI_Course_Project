magic
tech scmos
timestamp 1732011070
<< nwell >>
rect 3860 -1390 3884 -1366
rect 3899 -1376 3933 -1370
rect 3899 -1406 3961 -1376
rect 3927 -1412 3961 -1406
rect 3860 -1445 3884 -1421
rect -102 -1527 -78 -1503
rect -63 -1513 -29 -1507
rect -63 -1543 -1 -1513
rect -35 -1549 -1 -1543
rect -102 -1582 -78 -1558
rect 1596 -1663 1620 -1601
rect 1646 -1662 1670 -1600
rect 1696 -1662 1720 -1600
rect 1743 -1662 1767 -1600
rect 385 -1741 421 -1701
rect 427 -1748 451 -1708
rect -111 -1886 -87 -1862
rect -72 -1872 -38 -1866
rect -72 -1902 -10 -1872
rect 2065 -1884 2089 -1832
rect 2103 -1884 2127 -1832
rect 2147 -1884 2171 -1832
rect 2185 -1884 2209 -1832
rect 2231 -1882 2255 -1830
rect -44 -1908 -10 -1902
rect -111 -1941 -87 -1917
rect 387 -2091 423 -2051
rect 429 -2098 453 -2058
rect 3900 -2200 3924 -2176
rect 3939 -2186 3973 -2180
rect 3939 -2216 4001 -2186
rect -84 -2245 -60 -2221
rect 3967 -2222 4001 -2216
rect -45 -2231 -11 -2225
rect -45 -2261 17 -2231
rect 3900 -2255 3924 -2231
rect -17 -2267 17 -2261
rect -84 -2300 -60 -2276
rect 395 -2383 431 -2343
rect 437 -2390 461 -2350
rect -91 -2588 -67 -2564
rect -52 -2574 -18 -2568
rect -52 -2604 10 -2574
rect -24 -2610 10 -2604
rect -91 -2643 -67 -2619
rect 3840 -2630 3864 -2606
rect 3879 -2616 3913 -2610
rect 3879 -2646 3941 -2616
rect 3907 -2652 3941 -2646
rect 3840 -2685 3864 -2661
rect 383 -2749 419 -2709
rect 425 -2756 449 -2716
rect 3797 -3166 3821 -3142
rect 3836 -3152 3870 -3146
rect 3836 -3182 3898 -3152
rect 3864 -3188 3898 -3182
rect 3797 -3221 3821 -3197
<< ntransistor >>
rect 3871 -1404 3873 -1398
rect 3910 -1453 3912 -1441
rect 3920 -1453 3922 -1441
rect 3938 -1453 3940 -1441
rect 3948 -1453 3950 -1441
rect 3871 -1459 3873 -1453
rect -91 -1541 -89 -1535
rect -52 -1590 -50 -1578
rect -42 -1590 -40 -1578
rect -24 -1590 -22 -1578
rect -14 -1590 -12 -1578
rect -91 -1596 -89 -1590
rect 396 -1784 398 -1764
rect 407 -1784 409 -1764
rect 438 -1766 440 -1756
rect -100 -1900 -98 -1894
rect -61 -1949 -59 -1937
rect -51 -1949 -49 -1937
rect -33 -1949 -31 -1937
rect -23 -1949 -21 -1937
rect 1543 -1943 1545 -1843
rect 1571 -1943 1573 -1843
rect 1598 -1943 1600 -1843
rect 1637 -1943 1639 -1843
rect 1665 -1943 1667 -1843
rect 1692 -1943 1694 -1843
rect 1732 -1942 1734 -1842
rect 1760 -1942 1762 -1842
rect 1787 -1942 1789 -1842
rect 1823 -1942 1825 -1842
rect 2076 -1916 2078 -1896
rect 2114 -1916 2116 -1896
rect 2158 -1916 2160 -1896
rect 2196 -1916 2198 -1896
rect 2242 -1914 2244 -1894
rect -100 -1955 -98 -1949
rect 398 -2134 400 -2114
rect 409 -2134 411 -2114
rect 440 -2116 442 -2106
rect 3911 -2214 3913 -2208
rect -73 -2259 -71 -2253
rect 3950 -2263 3952 -2251
rect 3960 -2263 3962 -2251
rect 3978 -2263 3980 -2251
rect 3988 -2263 3990 -2251
rect 3911 -2269 3913 -2263
rect -34 -2308 -32 -2296
rect -24 -2308 -22 -2296
rect -6 -2308 -4 -2296
rect 4 -2308 6 -2296
rect -73 -2314 -71 -2308
rect 406 -2426 408 -2406
rect 417 -2426 419 -2406
rect 448 -2408 450 -2398
rect -80 -2602 -78 -2596
rect -41 -2651 -39 -2639
rect -31 -2651 -29 -2639
rect -13 -2651 -11 -2639
rect -3 -2651 -1 -2639
rect 3851 -2644 3853 -2638
rect -80 -2657 -78 -2651
rect 3890 -2693 3892 -2681
rect 3900 -2693 3902 -2681
rect 3918 -2693 3920 -2681
rect 3928 -2693 3930 -2681
rect 3851 -2699 3853 -2693
rect 394 -2792 396 -2772
rect 405 -2792 407 -2772
rect 436 -2774 438 -2764
rect 3808 -3180 3810 -3174
rect 3847 -3229 3849 -3217
rect 3857 -3229 3859 -3217
rect 3875 -3229 3877 -3217
rect 3885 -3229 3887 -3217
rect 3808 -3235 3810 -3229
<< ptransistor >>
rect 3871 -1384 3873 -1372
rect 3910 -1400 3912 -1376
rect 3920 -1400 3922 -1376
rect 3938 -1406 3940 -1382
rect 3948 -1406 3950 -1382
rect 3871 -1439 3873 -1427
rect -91 -1521 -89 -1509
rect -52 -1537 -50 -1513
rect -42 -1537 -40 -1513
rect -24 -1543 -22 -1519
rect -14 -1543 -12 -1519
rect -91 -1576 -89 -1564
rect 1607 -1657 1609 -1607
rect 1657 -1656 1659 -1606
rect 1707 -1656 1709 -1606
rect 1754 -1656 1756 -1606
rect 396 -1735 398 -1715
rect 407 -1735 409 -1715
rect 438 -1742 440 -1722
rect -100 -1880 -98 -1868
rect -61 -1896 -59 -1872
rect -51 -1896 -49 -1872
rect -33 -1902 -31 -1878
rect -23 -1902 -21 -1878
rect -100 -1935 -98 -1923
rect 2076 -1878 2078 -1838
rect 2114 -1878 2116 -1838
rect 2158 -1878 2160 -1838
rect 2196 -1878 2198 -1838
rect 2242 -1876 2244 -1836
rect 398 -2085 400 -2065
rect 409 -2085 411 -2065
rect 440 -2092 442 -2072
rect 3911 -2194 3913 -2182
rect 3950 -2210 3952 -2186
rect 3960 -2210 3962 -2186
rect 3978 -2216 3980 -2192
rect 3988 -2216 3990 -2192
rect -73 -2239 -71 -2227
rect -34 -2255 -32 -2231
rect -24 -2255 -22 -2231
rect -6 -2261 -4 -2237
rect 4 -2261 6 -2237
rect 3911 -2249 3913 -2237
rect -73 -2294 -71 -2282
rect 406 -2377 408 -2357
rect 417 -2377 419 -2357
rect 448 -2384 450 -2364
rect -80 -2582 -78 -2570
rect -41 -2598 -39 -2574
rect -31 -2598 -29 -2574
rect -13 -2604 -11 -2580
rect -3 -2604 -1 -2580
rect -80 -2637 -78 -2625
rect 3851 -2624 3853 -2612
rect 3890 -2640 3892 -2616
rect 3900 -2640 3902 -2616
rect 3918 -2646 3920 -2622
rect 3928 -2646 3930 -2622
rect 3851 -2679 3853 -2667
rect 394 -2743 396 -2723
rect 405 -2743 407 -2723
rect 436 -2750 438 -2730
rect 3808 -3160 3810 -3148
rect 3847 -3176 3849 -3152
rect 3857 -3176 3859 -3152
rect 3875 -3182 3877 -3158
rect 3885 -3182 3887 -3158
rect 3808 -3215 3810 -3203
<< ndiffusion >>
rect 3870 -1404 3871 -1398
rect 3873 -1404 3874 -1398
rect 3909 -1453 3910 -1441
rect 3912 -1453 3920 -1441
rect 3922 -1453 3923 -1441
rect 3937 -1453 3938 -1441
rect 3940 -1453 3948 -1441
rect 3950 -1453 3951 -1441
rect 3870 -1459 3871 -1453
rect 3873 -1459 3874 -1453
rect -92 -1541 -91 -1535
rect -89 -1541 -88 -1535
rect -53 -1590 -52 -1578
rect -50 -1590 -42 -1578
rect -40 -1590 -39 -1578
rect -25 -1590 -24 -1578
rect -22 -1590 -14 -1578
rect -12 -1590 -11 -1578
rect -92 -1596 -91 -1590
rect -89 -1596 -88 -1590
rect 395 -1784 396 -1764
rect 398 -1784 407 -1764
rect 409 -1784 410 -1764
rect 437 -1766 438 -1756
rect 440 -1766 441 -1756
rect -101 -1900 -100 -1894
rect -98 -1900 -97 -1894
rect -62 -1949 -61 -1937
rect -59 -1949 -51 -1937
rect -49 -1949 -48 -1937
rect -34 -1949 -33 -1937
rect -31 -1949 -23 -1937
rect -21 -1949 -20 -1937
rect 1542 -1943 1543 -1843
rect 1545 -1943 1546 -1843
rect 1570 -1943 1571 -1843
rect 1573 -1943 1574 -1843
rect 1597 -1943 1598 -1843
rect 1600 -1943 1601 -1843
rect 1636 -1943 1637 -1843
rect 1639 -1943 1640 -1843
rect 1664 -1943 1665 -1843
rect 1667 -1943 1668 -1843
rect 1691 -1943 1692 -1843
rect 1694 -1943 1695 -1843
rect 1731 -1942 1732 -1842
rect 1734 -1942 1735 -1842
rect 1759 -1942 1760 -1842
rect 1762 -1942 1763 -1842
rect 1786 -1942 1787 -1842
rect 1789 -1942 1790 -1842
rect 1822 -1942 1823 -1842
rect 1825 -1942 1826 -1842
rect 2075 -1916 2076 -1896
rect 2078 -1916 2079 -1896
rect 2113 -1916 2114 -1896
rect 2116 -1916 2117 -1896
rect 2157 -1916 2158 -1896
rect 2160 -1916 2161 -1896
rect 2195 -1916 2196 -1896
rect 2198 -1916 2199 -1896
rect 2241 -1914 2242 -1894
rect 2244 -1914 2245 -1894
rect -101 -1955 -100 -1949
rect -98 -1955 -97 -1949
rect 397 -2134 398 -2114
rect 400 -2134 409 -2114
rect 411 -2134 412 -2114
rect 439 -2116 440 -2106
rect 442 -2116 443 -2106
rect 3910 -2214 3911 -2208
rect 3913 -2214 3914 -2208
rect -74 -2259 -73 -2253
rect -71 -2259 -70 -2253
rect 3949 -2263 3950 -2251
rect 3952 -2263 3960 -2251
rect 3962 -2263 3963 -2251
rect 3977 -2263 3978 -2251
rect 3980 -2263 3988 -2251
rect 3990 -2263 3991 -2251
rect 3910 -2269 3911 -2263
rect 3913 -2269 3914 -2263
rect -35 -2308 -34 -2296
rect -32 -2308 -24 -2296
rect -22 -2308 -21 -2296
rect -7 -2308 -6 -2296
rect -4 -2308 4 -2296
rect 6 -2308 7 -2296
rect -74 -2314 -73 -2308
rect -71 -2314 -70 -2308
rect 405 -2426 406 -2406
rect 408 -2426 417 -2406
rect 419 -2426 420 -2406
rect 447 -2408 448 -2398
rect 450 -2408 451 -2398
rect -81 -2602 -80 -2596
rect -78 -2602 -77 -2596
rect -42 -2651 -41 -2639
rect -39 -2651 -31 -2639
rect -29 -2651 -28 -2639
rect -14 -2651 -13 -2639
rect -11 -2651 -3 -2639
rect -1 -2651 0 -2639
rect 3850 -2644 3851 -2638
rect 3853 -2644 3854 -2638
rect -81 -2657 -80 -2651
rect -78 -2657 -77 -2651
rect 3889 -2693 3890 -2681
rect 3892 -2693 3900 -2681
rect 3902 -2693 3903 -2681
rect 3917 -2693 3918 -2681
rect 3920 -2693 3928 -2681
rect 3930 -2693 3931 -2681
rect 3850 -2699 3851 -2693
rect 3853 -2699 3854 -2693
rect 393 -2792 394 -2772
rect 396 -2792 405 -2772
rect 407 -2792 408 -2772
rect 435 -2774 436 -2764
rect 438 -2774 439 -2764
rect 3807 -3180 3808 -3174
rect 3810 -3180 3811 -3174
rect 3846 -3229 3847 -3217
rect 3849 -3229 3857 -3217
rect 3859 -3229 3860 -3217
rect 3874 -3229 3875 -3217
rect 3877 -3229 3885 -3217
rect 3887 -3229 3888 -3217
rect 3807 -3235 3808 -3229
rect 3810 -3235 3811 -3229
<< pdiffusion >>
rect 3870 -1384 3871 -1372
rect 3873 -1384 3874 -1372
rect 3909 -1400 3910 -1376
rect 3912 -1400 3914 -1376
rect 3918 -1400 3920 -1376
rect 3922 -1400 3923 -1376
rect 3937 -1406 3938 -1382
rect 3940 -1406 3942 -1382
rect 3946 -1406 3948 -1382
rect 3950 -1406 3951 -1382
rect 3870 -1439 3871 -1427
rect 3873 -1439 3874 -1427
rect -92 -1521 -91 -1509
rect -89 -1521 -88 -1509
rect -53 -1537 -52 -1513
rect -50 -1537 -48 -1513
rect -44 -1537 -42 -1513
rect -40 -1537 -39 -1513
rect -25 -1543 -24 -1519
rect -22 -1543 -20 -1519
rect -16 -1543 -14 -1519
rect -12 -1543 -11 -1519
rect -92 -1576 -91 -1564
rect -89 -1576 -88 -1564
rect 1606 -1657 1607 -1607
rect 1609 -1657 1610 -1607
rect 1656 -1656 1657 -1606
rect 1659 -1656 1660 -1606
rect 1706 -1656 1707 -1606
rect 1709 -1656 1710 -1606
rect 1753 -1656 1754 -1606
rect 1756 -1656 1757 -1606
rect 395 -1735 396 -1715
rect 398 -1735 402 -1715
rect 406 -1735 407 -1715
rect 409 -1735 410 -1715
rect 437 -1742 438 -1722
rect 440 -1742 441 -1722
rect -101 -1880 -100 -1868
rect -98 -1880 -97 -1868
rect -62 -1896 -61 -1872
rect -59 -1896 -57 -1872
rect -53 -1896 -51 -1872
rect -49 -1896 -48 -1872
rect -34 -1902 -33 -1878
rect -31 -1902 -29 -1878
rect -25 -1902 -23 -1878
rect -21 -1902 -20 -1878
rect -101 -1935 -100 -1923
rect -98 -1935 -97 -1923
rect 2075 -1878 2076 -1838
rect 2078 -1878 2079 -1838
rect 2113 -1878 2114 -1838
rect 2116 -1878 2117 -1838
rect 2157 -1878 2158 -1838
rect 2160 -1878 2161 -1838
rect 2195 -1878 2196 -1838
rect 2198 -1878 2199 -1838
rect 2241 -1876 2242 -1836
rect 2244 -1876 2245 -1836
rect 397 -2085 398 -2065
rect 400 -2085 404 -2065
rect 408 -2085 409 -2065
rect 411 -2085 412 -2065
rect 439 -2092 440 -2072
rect 442 -2092 443 -2072
rect 3910 -2194 3911 -2182
rect 3913 -2194 3914 -2182
rect 3949 -2210 3950 -2186
rect 3952 -2210 3954 -2186
rect 3958 -2210 3960 -2186
rect 3962 -2210 3963 -2186
rect 3977 -2216 3978 -2192
rect 3980 -2216 3982 -2192
rect 3986 -2216 3988 -2192
rect 3990 -2216 3991 -2192
rect -74 -2239 -73 -2227
rect -71 -2239 -70 -2227
rect -35 -2255 -34 -2231
rect -32 -2255 -30 -2231
rect -26 -2255 -24 -2231
rect -22 -2255 -21 -2231
rect -7 -2261 -6 -2237
rect -4 -2261 -2 -2237
rect 2 -2261 4 -2237
rect 6 -2261 7 -2237
rect 3910 -2249 3911 -2237
rect 3913 -2249 3914 -2237
rect -74 -2294 -73 -2282
rect -71 -2294 -70 -2282
rect 405 -2377 406 -2357
rect 408 -2377 412 -2357
rect 416 -2377 417 -2357
rect 419 -2377 420 -2357
rect 447 -2384 448 -2364
rect 450 -2384 451 -2364
rect -81 -2582 -80 -2570
rect -78 -2582 -77 -2570
rect -42 -2598 -41 -2574
rect -39 -2598 -37 -2574
rect -33 -2598 -31 -2574
rect -29 -2598 -28 -2574
rect -14 -2604 -13 -2580
rect -11 -2604 -9 -2580
rect -5 -2604 -3 -2580
rect -1 -2604 0 -2580
rect -81 -2637 -80 -2625
rect -78 -2637 -77 -2625
rect 3850 -2624 3851 -2612
rect 3853 -2624 3854 -2612
rect 3889 -2640 3890 -2616
rect 3892 -2640 3894 -2616
rect 3898 -2640 3900 -2616
rect 3902 -2640 3903 -2616
rect 3917 -2646 3918 -2622
rect 3920 -2646 3922 -2622
rect 3926 -2646 3928 -2622
rect 3930 -2646 3931 -2622
rect 3850 -2679 3851 -2667
rect 3853 -2679 3854 -2667
rect 393 -2743 394 -2723
rect 396 -2743 400 -2723
rect 404 -2743 405 -2723
rect 407 -2743 408 -2723
rect 435 -2750 436 -2730
rect 438 -2750 439 -2730
rect 3807 -3160 3808 -3148
rect 3810 -3160 3811 -3148
rect 3846 -3176 3847 -3152
rect 3849 -3176 3851 -3152
rect 3855 -3176 3857 -3152
rect 3859 -3176 3860 -3152
rect 3874 -3182 3875 -3158
rect 3877 -3182 3879 -3158
rect 3883 -3182 3885 -3158
rect 3887 -3182 3888 -3158
rect 3807 -3215 3808 -3203
rect 3810 -3215 3811 -3203
<< ndcontact >>
rect 3866 -1404 3870 -1398
rect 3874 -1404 3878 -1398
rect 3905 -1453 3909 -1441
rect 3923 -1453 3927 -1441
rect 3933 -1453 3937 -1441
rect 3951 -1453 3955 -1441
rect 3866 -1459 3870 -1453
rect 3874 -1459 3878 -1453
rect -96 -1541 -92 -1535
rect -88 -1541 -84 -1535
rect -57 -1590 -53 -1578
rect -39 -1590 -35 -1578
rect -29 -1590 -25 -1578
rect -11 -1590 -7 -1578
rect -96 -1596 -92 -1590
rect -88 -1596 -84 -1590
rect 391 -1784 395 -1764
rect 410 -1784 414 -1764
rect 433 -1766 437 -1756
rect 441 -1766 445 -1756
rect -105 -1900 -101 -1894
rect -97 -1900 -93 -1894
rect -66 -1949 -62 -1937
rect -48 -1949 -44 -1937
rect -38 -1949 -34 -1937
rect -20 -1949 -16 -1937
rect 1538 -1943 1542 -1843
rect 1546 -1943 1550 -1843
rect 1566 -1943 1570 -1843
rect 1574 -1943 1578 -1843
rect 1593 -1943 1597 -1843
rect 1601 -1943 1605 -1843
rect 1632 -1943 1636 -1843
rect 1640 -1943 1644 -1843
rect 1660 -1943 1664 -1843
rect 1668 -1943 1672 -1843
rect 1687 -1943 1691 -1843
rect 1695 -1943 1699 -1843
rect 1727 -1942 1731 -1842
rect 1735 -1942 1739 -1842
rect 1755 -1942 1759 -1842
rect 1763 -1942 1767 -1842
rect 1782 -1942 1786 -1842
rect 1790 -1942 1794 -1842
rect 1818 -1942 1822 -1842
rect 1826 -1942 1830 -1842
rect 2071 -1916 2075 -1896
rect 2079 -1916 2083 -1896
rect 2109 -1916 2113 -1896
rect 2117 -1916 2121 -1896
rect 2153 -1916 2157 -1896
rect 2161 -1916 2165 -1896
rect 2191 -1916 2195 -1896
rect 2199 -1916 2203 -1896
rect 2237 -1914 2241 -1894
rect 2245 -1914 2249 -1894
rect -105 -1955 -101 -1949
rect -97 -1955 -93 -1949
rect 393 -2134 397 -2114
rect 412 -2134 416 -2114
rect 435 -2116 439 -2106
rect 443 -2116 447 -2106
rect 3906 -2214 3910 -2208
rect 3914 -2214 3918 -2208
rect -78 -2259 -74 -2253
rect -70 -2259 -66 -2253
rect 3945 -2263 3949 -2251
rect 3963 -2263 3967 -2251
rect 3973 -2263 3977 -2251
rect 3991 -2263 3995 -2251
rect 3906 -2269 3910 -2263
rect 3914 -2269 3918 -2263
rect -39 -2308 -35 -2296
rect -21 -2308 -17 -2296
rect -11 -2308 -7 -2296
rect 7 -2308 11 -2296
rect -78 -2314 -74 -2308
rect -70 -2314 -66 -2308
rect 401 -2426 405 -2406
rect 420 -2426 424 -2406
rect 443 -2408 447 -2398
rect 451 -2408 455 -2398
rect -85 -2602 -81 -2596
rect -77 -2602 -73 -2596
rect -46 -2651 -42 -2639
rect -28 -2651 -24 -2639
rect -18 -2651 -14 -2639
rect 0 -2651 4 -2639
rect 3846 -2644 3850 -2638
rect 3854 -2644 3858 -2638
rect -85 -2657 -81 -2651
rect -77 -2657 -73 -2651
rect 3885 -2693 3889 -2681
rect 3903 -2693 3907 -2681
rect 3913 -2693 3917 -2681
rect 3931 -2693 3935 -2681
rect 3846 -2699 3850 -2693
rect 3854 -2699 3858 -2693
rect 389 -2792 393 -2772
rect 408 -2792 412 -2772
rect 431 -2774 435 -2764
rect 439 -2774 443 -2764
rect 3803 -3180 3807 -3174
rect 3811 -3180 3815 -3174
rect 3842 -3229 3846 -3217
rect 3860 -3229 3864 -3217
rect 3870 -3229 3874 -3217
rect 3888 -3229 3892 -3217
rect 3803 -3235 3807 -3229
rect 3811 -3235 3815 -3229
<< pdcontact >>
rect 3866 -1384 3870 -1372
rect 3874 -1384 3878 -1372
rect 3905 -1400 3909 -1376
rect 3914 -1400 3918 -1376
rect 3923 -1400 3927 -1376
rect 3933 -1406 3937 -1382
rect 3942 -1406 3946 -1382
rect 3951 -1406 3955 -1382
rect 3866 -1439 3870 -1427
rect 3874 -1439 3878 -1427
rect -96 -1521 -92 -1509
rect -88 -1521 -84 -1509
rect -57 -1537 -53 -1513
rect -48 -1537 -44 -1513
rect -39 -1537 -35 -1513
rect -29 -1543 -25 -1519
rect -20 -1543 -16 -1519
rect -11 -1543 -7 -1519
rect -96 -1576 -92 -1564
rect -88 -1576 -84 -1564
rect 1602 -1657 1606 -1607
rect 1610 -1657 1614 -1607
rect 1652 -1656 1656 -1606
rect 1660 -1656 1664 -1606
rect 1702 -1656 1706 -1606
rect 1710 -1656 1714 -1606
rect 1749 -1656 1753 -1606
rect 1757 -1656 1761 -1606
rect 391 -1735 395 -1715
rect 402 -1735 406 -1715
rect 410 -1735 414 -1715
rect 433 -1742 437 -1722
rect 441 -1742 445 -1722
rect -105 -1880 -101 -1868
rect -97 -1880 -93 -1868
rect -66 -1896 -62 -1872
rect -57 -1896 -53 -1872
rect -48 -1896 -44 -1872
rect -38 -1902 -34 -1878
rect -29 -1902 -25 -1878
rect -20 -1902 -16 -1878
rect -105 -1935 -101 -1923
rect -97 -1935 -93 -1923
rect 2071 -1878 2075 -1838
rect 2079 -1878 2083 -1838
rect 2109 -1878 2113 -1838
rect 2117 -1878 2121 -1838
rect 2153 -1878 2157 -1838
rect 2161 -1878 2165 -1838
rect 2191 -1878 2195 -1838
rect 2199 -1878 2203 -1838
rect 2237 -1876 2241 -1836
rect 2245 -1876 2249 -1836
rect 393 -2085 397 -2065
rect 404 -2085 408 -2065
rect 412 -2085 416 -2065
rect 435 -2092 439 -2072
rect 443 -2092 447 -2072
rect 3906 -2194 3910 -2182
rect 3914 -2194 3918 -2182
rect 3945 -2210 3949 -2186
rect 3954 -2210 3958 -2186
rect 3963 -2210 3967 -2186
rect 3973 -2216 3977 -2192
rect 3982 -2216 3986 -2192
rect 3991 -2216 3995 -2192
rect -78 -2239 -74 -2227
rect -70 -2239 -66 -2227
rect -39 -2255 -35 -2231
rect -30 -2255 -26 -2231
rect -21 -2255 -17 -2231
rect -11 -2261 -7 -2237
rect -2 -2261 2 -2237
rect 7 -2261 11 -2237
rect 3906 -2249 3910 -2237
rect 3914 -2249 3918 -2237
rect -78 -2294 -74 -2282
rect -70 -2294 -66 -2282
rect 401 -2377 405 -2357
rect 412 -2377 416 -2357
rect 420 -2377 424 -2357
rect 443 -2384 447 -2364
rect 451 -2384 455 -2364
rect -85 -2582 -81 -2570
rect -77 -2582 -73 -2570
rect -46 -2598 -42 -2574
rect -37 -2598 -33 -2574
rect -28 -2598 -24 -2574
rect -18 -2604 -14 -2580
rect -9 -2604 -5 -2580
rect 0 -2604 4 -2580
rect -85 -2637 -81 -2625
rect -77 -2637 -73 -2625
rect 3846 -2624 3850 -2612
rect 3854 -2624 3858 -2612
rect 3885 -2640 3889 -2616
rect 3894 -2640 3898 -2616
rect 3903 -2640 3907 -2616
rect 3913 -2646 3917 -2622
rect 3922 -2646 3926 -2622
rect 3931 -2646 3935 -2622
rect 3846 -2679 3850 -2667
rect 3854 -2679 3858 -2667
rect 389 -2743 393 -2723
rect 400 -2743 404 -2723
rect 408 -2743 412 -2723
rect 431 -2750 435 -2730
rect 439 -2750 443 -2730
rect 3803 -3160 3807 -3148
rect 3811 -3160 3815 -3148
rect 3842 -3176 3846 -3152
rect 3851 -3176 3855 -3152
rect 3860 -3176 3864 -3152
rect 3870 -3182 3874 -3158
rect 3879 -3182 3883 -3158
rect 3888 -3182 3892 -3158
rect 3803 -3215 3807 -3203
rect 3811 -3215 3815 -3203
<< psubstratepcontact >>
rect 447 -1775 452 -1771
rect 449 -2125 454 -2121
rect 457 -2417 462 -2413
rect 445 -2783 450 -2779
<< nsubstratencontact >>
rect 1597 -1601 1601 -1596
rect 1647 -1600 1651 -1595
rect 1697 -1600 1701 -1595
rect 1744 -1600 1748 -1595
rect 391 -1710 395 -1704
rect 443 -1715 447 -1711
rect 2066 -1832 2070 -1828
rect 2104 -1832 2108 -1828
rect 2148 -1832 2152 -1828
rect 2186 -1832 2190 -1828
rect 2232 -1830 2236 -1826
rect 393 -2060 397 -2054
rect 445 -2065 449 -2061
rect 401 -2352 405 -2346
rect 453 -2357 457 -2353
rect 389 -2718 393 -2712
rect 441 -2723 445 -2719
<< polysilicon >>
rect 3871 -1372 3873 -1369
rect 3910 -1376 3912 -1373
rect 3920 -1376 3922 -1373
rect 3871 -1398 3873 -1384
rect 3938 -1382 3940 -1379
rect 3948 -1382 3950 -1379
rect 3871 -1407 3873 -1404
rect 3910 -1409 3912 -1400
rect 3920 -1410 3922 -1400
rect 3871 -1427 3873 -1424
rect 3871 -1453 3873 -1439
rect 3910 -1441 3912 -1414
rect 3920 -1441 3922 -1415
rect 3938 -1417 3940 -1406
rect 3938 -1441 3940 -1421
rect 3948 -1428 3950 -1406
rect 3948 -1441 3950 -1432
rect 3910 -1456 3912 -1453
rect 3920 -1456 3922 -1453
rect 3938 -1456 3940 -1453
rect 3948 -1456 3950 -1453
rect 3871 -1462 3873 -1459
rect -91 -1509 -89 -1506
rect -52 -1513 -50 -1510
rect -42 -1513 -40 -1510
rect -91 -1535 -89 -1521
rect -24 -1519 -22 -1516
rect -14 -1519 -12 -1516
rect -91 -1544 -89 -1541
rect -52 -1546 -50 -1537
rect -42 -1547 -40 -1537
rect -91 -1564 -89 -1561
rect -91 -1590 -89 -1576
rect -52 -1578 -50 -1551
rect -42 -1578 -40 -1552
rect -24 -1554 -22 -1543
rect -24 -1578 -22 -1558
rect -14 -1565 -12 -1543
rect -14 -1578 -12 -1569
rect -52 -1593 -50 -1590
rect -42 -1593 -40 -1590
rect -24 -1593 -22 -1590
rect -14 -1593 -12 -1590
rect -91 -1599 -89 -1596
rect 1607 -1607 1609 -1604
rect 1657 -1606 1659 -1603
rect 1707 -1606 1709 -1603
rect 1754 -1606 1756 -1603
rect 1607 -1680 1609 -1657
rect 1657 -1679 1659 -1656
rect 1707 -1679 1709 -1656
rect 1754 -1679 1756 -1656
rect 396 -1715 398 -1712
rect 407 -1715 409 -1712
rect 438 -1722 440 -1718
rect 396 -1764 398 -1735
rect 407 -1764 409 -1735
rect 438 -1756 440 -1742
rect 438 -1769 440 -1766
rect 396 -1787 398 -1784
rect 407 -1787 409 -1784
rect 2076 -1838 2078 -1835
rect 2114 -1838 2116 -1835
rect 2158 -1838 2160 -1835
rect 2196 -1838 2198 -1835
rect 2242 -1836 2244 -1833
rect 1543 -1843 1545 -1840
rect 1571 -1843 1573 -1840
rect 1598 -1843 1600 -1840
rect 1637 -1843 1639 -1840
rect 1665 -1843 1667 -1840
rect 1692 -1843 1694 -1840
rect 1732 -1842 1734 -1839
rect 1760 -1842 1762 -1839
rect 1787 -1842 1789 -1839
rect 1823 -1842 1825 -1839
rect -100 -1868 -98 -1865
rect -61 -1872 -59 -1869
rect -51 -1872 -49 -1869
rect -100 -1894 -98 -1880
rect -33 -1878 -31 -1875
rect -23 -1878 -21 -1875
rect -100 -1903 -98 -1900
rect -61 -1905 -59 -1896
rect -51 -1906 -49 -1896
rect -100 -1923 -98 -1920
rect -100 -1949 -98 -1935
rect -61 -1937 -59 -1910
rect -51 -1937 -49 -1911
rect -33 -1913 -31 -1902
rect -33 -1937 -31 -1917
rect -23 -1924 -21 -1902
rect -23 -1937 -21 -1928
rect 2076 -1896 2078 -1878
rect 2114 -1896 2116 -1878
rect 2158 -1896 2160 -1878
rect 2196 -1896 2198 -1878
rect 2242 -1894 2244 -1876
rect 2076 -1920 2078 -1916
rect 2114 -1920 2116 -1916
rect 2158 -1920 2160 -1916
rect 2196 -1920 2198 -1916
rect 2242 -1918 2244 -1914
rect -61 -1952 -59 -1949
rect -51 -1952 -49 -1949
rect -33 -1952 -31 -1949
rect -23 -1952 -21 -1949
rect 1543 -1955 1545 -1943
rect 1571 -1955 1573 -1943
rect 1598 -1955 1600 -1943
rect 1637 -1955 1639 -1943
rect 1665 -1955 1667 -1943
rect 1692 -1955 1694 -1943
rect 1732 -1954 1734 -1942
rect 1760 -1954 1762 -1942
rect 1787 -1954 1789 -1942
rect 1823 -1954 1825 -1942
rect -100 -1958 -98 -1955
rect 398 -2065 400 -2062
rect 409 -2065 411 -2062
rect 440 -2072 442 -2068
rect 398 -2114 400 -2085
rect 409 -2114 411 -2085
rect 440 -2106 442 -2092
rect 440 -2119 442 -2116
rect 398 -2137 400 -2134
rect 409 -2137 411 -2134
rect 3911 -2182 3913 -2179
rect 3950 -2186 3952 -2183
rect 3960 -2186 3962 -2183
rect 3911 -2208 3913 -2194
rect 3978 -2192 3980 -2189
rect 3988 -2192 3990 -2189
rect 3911 -2217 3913 -2214
rect 3950 -2219 3952 -2210
rect 3960 -2220 3962 -2210
rect -73 -2227 -71 -2224
rect -34 -2231 -32 -2228
rect -24 -2231 -22 -2228
rect -73 -2253 -71 -2239
rect -6 -2237 -4 -2234
rect 4 -2237 6 -2234
rect 3911 -2237 3913 -2234
rect -73 -2262 -71 -2259
rect -34 -2264 -32 -2255
rect -24 -2265 -22 -2255
rect -73 -2282 -71 -2279
rect -73 -2308 -71 -2294
rect -34 -2296 -32 -2269
rect -24 -2296 -22 -2270
rect -6 -2272 -4 -2261
rect -6 -2296 -4 -2276
rect 4 -2283 6 -2261
rect 3911 -2263 3913 -2249
rect 3950 -2251 3952 -2224
rect 3960 -2251 3962 -2225
rect 3978 -2227 3980 -2216
rect 3978 -2251 3980 -2231
rect 3988 -2238 3990 -2216
rect 3988 -2251 3990 -2242
rect 3950 -2266 3952 -2263
rect 3960 -2266 3962 -2263
rect 3978 -2266 3980 -2263
rect 3988 -2266 3990 -2263
rect 3911 -2272 3913 -2269
rect 4 -2296 6 -2287
rect -34 -2311 -32 -2308
rect -24 -2311 -22 -2308
rect -6 -2311 -4 -2308
rect 4 -2311 6 -2308
rect -73 -2317 -71 -2314
rect 406 -2357 408 -2354
rect 417 -2357 419 -2354
rect 448 -2364 450 -2360
rect 406 -2406 408 -2377
rect 417 -2406 419 -2377
rect 448 -2398 450 -2384
rect 448 -2411 450 -2408
rect 406 -2429 408 -2426
rect 417 -2429 419 -2426
rect -80 -2570 -78 -2567
rect -41 -2574 -39 -2571
rect -31 -2574 -29 -2571
rect -80 -2596 -78 -2582
rect -13 -2580 -11 -2577
rect -3 -2580 -1 -2577
rect -80 -2605 -78 -2602
rect -41 -2607 -39 -2598
rect -31 -2608 -29 -2598
rect -80 -2625 -78 -2622
rect -80 -2651 -78 -2637
rect -41 -2639 -39 -2612
rect -31 -2639 -29 -2613
rect -13 -2615 -11 -2604
rect -13 -2639 -11 -2619
rect -3 -2626 -1 -2604
rect 3851 -2612 3853 -2609
rect 3890 -2616 3892 -2613
rect 3900 -2616 3902 -2613
rect -3 -2639 -1 -2630
rect 3851 -2638 3853 -2624
rect 3918 -2622 3920 -2619
rect 3928 -2622 3930 -2619
rect 3851 -2647 3853 -2644
rect 3890 -2649 3892 -2640
rect -41 -2654 -39 -2651
rect -31 -2654 -29 -2651
rect -13 -2654 -11 -2651
rect -3 -2654 -1 -2651
rect 3900 -2650 3902 -2640
rect -80 -2660 -78 -2657
rect 3851 -2667 3853 -2664
rect 3851 -2693 3853 -2679
rect 3890 -2681 3892 -2654
rect 3900 -2681 3902 -2655
rect 3918 -2657 3920 -2646
rect 3918 -2681 3920 -2661
rect 3928 -2668 3930 -2646
rect 3928 -2681 3930 -2672
rect 3890 -2696 3892 -2693
rect 3900 -2696 3902 -2693
rect 3918 -2696 3920 -2693
rect 3928 -2696 3930 -2693
rect 3851 -2702 3853 -2699
rect 394 -2723 396 -2720
rect 405 -2723 407 -2720
rect 436 -2730 438 -2726
rect 394 -2772 396 -2743
rect 405 -2772 407 -2743
rect 436 -2764 438 -2750
rect 436 -2777 438 -2774
rect 394 -2795 396 -2792
rect 405 -2795 407 -2792
rect 3808 -3148 3810 -3145
rect 3847 -3152 3849 -3149
rect 3857 -3152 3859 -3149
rect 3808 -3174 3810 -3160
rect 3875 -3158 3877 -3155
rect 3885 -3158 3887 -3155
rect 3808 -3183 3810 -3180
rect 3847 -3185 3849 -3176
rect 3857 -3186 3859 -3176
rect 3808 -3203 3810 -3200
rect 3808 -3229 3810 -3215
rect 3847 -3217 3849 -3190
rect 3857 -3217 3859 -3191
rect 3875 -3193 3877 -3182
rect 3875 -3217 3877 -3197
rect 3885 -3204 3887 -3182
rect 3885 -3217 3887 -3208
rect 3847 -3232 3849 -3229
rect 3857 -3232 3859 -3229
rect 3875 -3232 3877 -3229
rect 3885 -3232 3887 -3229
rect 3808 -3238 3810 -3235
<< polycontact >>
rect 3867 -1395 3871 -1391
rect 3867 -1450 3871 -1446
rect 3936 -1421 3940 -1417
rect 3947 -1432 3951 -1428
rect -95 -1532 -91 -1528
rect -95 -1587 -91 -1583
rect -26 -1558 -22 -1554
rect -15 -1569 -11 -1565
rect 392 -1761 396 -1757
rect 403 -1754 407 -1750
rect 434 -1753 438 -1749
rect -104 -1891 -100 -1887
rect -104 -1946 -100 -1942
rect -35 -1917 -31 -1913
rect -24 -1928 -20 -1924
rect 394 -2111 398 -2107
rect 405 -2104 409 -2100
rect 436 -2103 440 -2099
rect 3907 -2205 3911 -2201
rect -77 -2250 -73 -2246
rect 3907 -2260 3911 -2256
rect -77 -2305 -73 -2301
rect -8 -2276 -4 -2272
rect 3976 -2231 3980 -2227
rect 3987 -2242 3991 -2238
rect 3 -2287 7 -2283
rect 402 -2403 406 -2399
rect 413 -2396 417 -2392
rect 444 -2395 448 -2391
rect -84 -2593 -80 -2589
rect -84 -2648 -80 -2644
rect -15 -2619 -11 -2615
rect -4 -2630 0 -2626
rect 3847 -2635 3851 -2631
rect 3847 -2690 3851 -2686
rect 3916 -2661 3920 -2657
rect 3927 -2672 3931 -2668
rect 390 -2769 394 -2765
rect 401 -2762 405 -2758
rect 432 -2761 436 -2757
rect 3804 -3171 3808 -3167
rect 3804 -3226 3808 -3222
rect 3873 -3197 3877 -3193
rect 3884 -3208 3888 -3204
<< metal1 >>
rect 3865 -1366 3893 -1363
rect 3866 -1372 3869 -1366
rect 3890 -1367 3893 -1366
rect 3890 -1370 3961 -1367
rect 3849 -1396 3852 -1393
rect 3857 -1395 3867 -1392
rect 3875 -1392 3878 -1384
rect 3905 -1376 3908 -1370
rect 3924 -1376 3927 -1370
rect 3875 -1395 3896 -1392
rect 3875 -1398 3878 -1395
rect 3866 -1408 3869 -1404
rect 3860 -1410 3884 -1408
rect 3860 -1411 3878 -1410
rect 3883 -1411 3884 -1410
rect 3893 -1418 3896 -1395
rect 3934 -1376 3954 -1373
rect 3934 -1382 3937 -1376
rect 3951 -1382 3954 -1376
rect 3915 -1403 3918 -1400
rect 3915 -1406 3933 -1403
rect 3943 -1413 3946 -1406
rect 3943 -1416 3960 -1413
rect 3865 -1419 3884 -1418
rect 3860 -1421 3884 -1419
rect 3893 -1421 3936 -1418
rect 3866 -1427 3869 -1421
rect 3957 -1427 3960 -1416
rect 3922 -1432 3947 -1429
rect 3957 -1431 3970 -1427
rect 3922 -1434 3925 -1432
rect 3849 -1450 3852 -1447
rect 3857 -1450 3867 -1447
rect 3875 -1447 3878 -1439
rect 3887 -1437 3925 -1434
rect 3957 -1435 3960 -1431
rect 3887 -1447 3890 -1437
rect 3928 -1438 3960 -1435
rect 3928 -1441 3931 -1438
rect 3875 -1450 3890 -1447
rect 3875 -1453 3878 -1450
rect 3927 -1444 3933 -1441
rect 3866 -1463 3869 -1459
rect 3887 -1460 3892 -1457
rect 3905 -1457 3908 -1453
rect 3952 -1457 3955 -1453
rect 3897 -1460 3961 -1457
rect 3887 -1463 3890 -1460
rect 3860 -1466 3890 -1463
rect 3966 -1471 3970 -1431
rect -97 -1503 -69 -1500
rect -96 -1509 -93 -1503
rect -72 -1504 -69 -1503
rect -72 -1507 -1 -1504
rect -113 -1533 -110 -1530
rect -105 -1532 -95 -1529
rect -87 -1529 -84 -1521
rect -57 -1513 -54 -1507
rect -38 -1513 -35 -1507
rect -87 -1532 -66 -1529
rect -87 -1535 -84 -1532
rect -96 -1545 -93 -1541
rect -102 -1547 -78 -1545
rect -102 -1548 -84 -1547
rect -79 -1548 -78 -1547
rect -69 -1555 -66 -1532
rect -28 -1513 -8 -1510
rect -28 -1519 -25 -1513
rect -11 -1519 -8 -1513
rect -47 -1540 -44 -1537
rect -47 -1543 -29 -1540
rect -19 -1550 -16 -1543
rect -19 -1553 -2 -1550
rect -97 -1556 -78 -1555
rect -102 -1558 -78 -1556
rect -69 -1558 -26 -1555
rect -96 -1564 -93 -1558
rect -5 -1564 -2 -1553
rect -40 -1569 -15 -1566
rect -5 -1568 8 -1564
rect -40 -1571 -37 -1569
rect -113 -1587 -110 -1584
rect -105 -1587 -95 -1584
rect -87 -1584 -84 -1576
rect -75 -1574 -37 -1571
rect -5 -1572 -2 -1568
rect -75 -1584 -72 -1574
rect -34 -1575 -2 -1572
rect -34 -1578 -31 -1575
rect -87 -1587 -72 -1584
rect -87 -1590 -84 -1587
rect -35 -1581 -29 -1578
rect -96 -1600 -93 -1596
rect -75 -1597 -70 -1594
rect -57 -1594 -54 -1590
rect -10 -1594 -7 -1590
rect -65 -1597 -1 -1594
rect -75 -1600 -72 -1597
rect -102 -1603 -72 -1600
rect 4 -1608 8 -1568
rect 1602 -1596 1606 -1587
rect 1652 -1595 1656 -1586
rect 1702 -1595 1706 -1586
rect 1749 -1595 1753 -1586
rect 1596 -1601 1597 -1596
rect 1601 -1601 1620 -1596
rect 1646 -1600 1647 -1595
rect 1651 -1600 1670 -1595
rect 1696 -1600 1697 -1595
rect 1701 -1600 1720 -1595
rect 1743 -1600 1744 -1595
rect 1748 -1600 1767 -1595
rect 1602 -1607 1606 -1601
rect 1652 -1606 1656 -1600
rect 1702 -1606 1706 -1600
rect 1749 -1606 1753 -1600
rect 1610 -1671 1614 -1657
rect 1660 -1670 1664 -1656
rect 1710 -1670 1714 -1656
rect 1757 -1670 1761 -1656
rect 391 -1704 414 -1700
rect 395 -1706 414 -1704
rect 391 -1715 395 -1710
rect 410 -1715 414 -1706
rect 427 -1711 451 -1710
rect 427 -1715 443 -1711
rect 447 -1715 451 -1711
rect 427 -1717 451 -1715
rect 433 -1722 437 -1717
rect 402 -1743 406 -1735
rect 402 -1747 414 -1743
rect 410 -1749 414 -1747
rect 441 -1749 445 -1742
rect 385 -1754 403 -1750
rect 410 -1753 434 -1749
rect 441 -1753 451 -1749
rect 385 -1761 392 -1757
rect 410 -1764 414 -1753
rect 441 -1756 445 -1753
rect 433 -1770 437 -1766
rect 427 -1771 452 -1770
rect 427 -1775 447 -1771
rect 427 -1776 452 -1775
rect 391 -1788 395 -1784
rect 391 -1792 407 -1788
rect 2071 -1825 2091 -1821
rect 2102 -1825 2133 -1821
rect 2145 -1825 2173 -1821
rect 2183 -1825 2204 -1821
rect 2220 -1823 2250 -1819
rect 2071 -1828 2075 -1825
rect 2109 -1828 2113 -1825
rect 2153 -1828 2157 -1825
rect 2191 -1828 2195 -1825
rect 2237 -1826 2241 -1823
rect 2065 -1832 2066 -1828
rect 2070 -1832 2075 -1828
rect 2103 -1832 2104 -1828
rect 2108 -1832 2113 -1828
rect 2147 -1832 2148 -1828
rect 2152 -1832 2157 -1828
rect 2185 -1832 2186 -1828
rect 2190 -1832 2195 -1828
rect 2231 -1830 2232 -1826
rect 2236 -1830 2241 -1826
rect 1538 -1843 1542 -1835
rect 1566 -1843 1570 -1835
rect 1593 -1843 1597 -1835
rect 1632 -1843 1636 -1835
rect 1660 -1843 1664 -1835
rect 1687 -1843 1691 -1835
rect 1727 -1842 1731 -1834
rect 1755 -1842 1759 -1834
rect 1782 -1842 1786 -1834
rect 1818 -1842 1822 -1834
rect 2071 -1838 2075 -1832
rect 2109 -1838 2113 -1832
rect 2153 -1838 2157 -1832
rect 2191 -1838 2195 -1832
rect 2237 -1836 2241 -1830
rect -106 -1862 -78 -1859
rect -105 -1868 -102 -1862
rect -81 -1863 -78 -1862
rect -81 -1866 -10 -1863
rect -122 -1892 -119 -1889
rect -114 -1891 -104 -1888
rect -96 -1888 -93 -1880
rect -66 -1872 -63 -1866
rect -47 -1872 -44 -1866
rect -96 -1891 -75 -1888
rect -96 -1894 -93 -1891
rect -105 -1904 -102 -1900
rect -111 -1906 -87 -1904
rect -111 -1907 -93 -1906
rect -88 -1907 -87 -1906
rect -78 -1914 -75 -1891
rect -37 -1872 -17 -1869
rect -37 -1878 -34 -1872
rect -20 -1878 -17 -1872
rect -56 -1899 -53 -1896
rect -56 -1902 -38 -1899
rect -28 -1909 -25 -1902
rect -28 -1912 -11 -1909
rect -106 -1915 -87 -1914
rect -111 -1917 -87 -1915
rect -78 -1917 -35 -1914
rect -105 -1923 -102 -1917
rect -14 -1923 -11 -1912
rect -49 -1928 -24 -1925
rect -14 -1927 -1 -1923
rect -49 -1930 -46 -1928
rect -122 -1946 -119 -1943
rect -114 -1946 -104 -1943
rect -96 -1943 -93 -1935
rect -84 -1933 -46 -1930
rect -14 -1931 -11 -1927
rect -84 -1943 -81 -1933
rect -43 -1934 -11 -1931
rect -43 -1937 -40 -1934
rect -96 -1946 -81 -1943
rect -96 -1949 -93 -1946
rect -44 -1940 -38 -1937
rect -105 -1959 -102 -1955
rect -84 -1956 -79 -1953
rect -66 -1953 -63 -1949
rect -19 -1953 -16 -1949
rect -74 -1956 -10 -1953
rect -84 -1959 -81 -1956
rect -111 -1962 -81 -1959
rect -5 -1967 -1 -1927
rect 2079 -1896 2083 -1878
rect 2117 -1896 2121 -1878
rect 2161 -1896 2165 -1878
rect 2199 -1896 2203 -1878
rect 2245 -1894 2249 -1876
rect 2071 -1925 2075 -1916
rect 2109 -1925 2113 -1916
rect 2153 -1925 2157 -1916
rect 2191 -1925 2195 -1916
rect 2237 -1923 2241 -1914
rect 2071 -1929 2091 -1925
rect 2102 -1929 2133 -1925
rect 2145 -1929 2173 -1925
rect 2183 -1929 2200 -1925
rect 2220 -1927 2246 -1923
rect 1546 -1949 1550 -1943
rect 1574 -1949 1578 -1943
rect 1601 -1949 1605 -1943
rect 1640 -1949 1644 -1943
rect 1668 -1949 1672 -1943
rect 1695 -1949 1699 -1943
rect 1735 -1948 1739 -1942
rect 1763 -1948 1767 -1942
rect 1790 -1948 1794 -1942
rect 1826 -1948 1830 -1942
rect 393 -2054 416 -2050
rect 397 -2056 416 -2054
rect 393 -2065 397 -2060
rect 412 -2065 416 -2056
rect 429 -2061 453 -2060
rect 429 -2065 445 -2061
rect 449 -2065 453 -2061
rect 429 -2067 453 -2065
rect 435 -2072 439 -2067
rect 404 -2093 408 -2085
rect 404 -2097 416 -2093
rect 412 -2099 416 -2097
rect 443 -2099 447 -2092
rect 387 -2104 405 -2100
rect 412 -2103 436 -2099
rect 443 -2103 453 -2099
rect 387 -2111 394 -2107
rect 412 -2114 416 -2103
rect 443 -2106 447 -2103
rect 435 -2120 439 -2116
rect 429 -2121 454 -2120
rect 429 -2125 449 -2121
rect 429 -2126 454 -2125
rect 393 -2138 397 -2134
rect 393 -2142 409 -2138
rect 3905 -2176 3933 -2173
rect 3906 -2182 3909 -2176
rect 3930 -2177 3933 -2176
rect 3930 -2180 4001 -2177
rect 3889 -2206 3892 -2203
rect 3897 -2205 3907 -2202
rect 3915 -2202 3918 -2194
rect 3945 -2186 3948 -2180
rect 3964 -2186 3967 -2180
rect 3915 -2205 3936 -2202
rect 3915 -2208 3918 -2205
rect 3906 -2218 3909 -2214
rect -79 -2221 -51 -2218
rect 3900 -2220 3924 -2218
rect 3900 -2221 3918 -2220
rect -78 -2227 -75 -2221
rect -54 -2222 -51 -2221
rect -54 -2225 17 -2222
rect -95 -2251 -92 -2248
rect -87 -2250 -77 -2247
rect -69 -2247 -66 -2239
rect -39 -2231 -36 -2225
rect -20 -2231 -17 -2225
rect -69 -2250 -48 -2247
rect -69 -2253 -66 -2250
rect -78 -2263 -75 -2259
rect -84 -2265 -60 -2263
rect -84 -2266 -66 -2265
rect -61 -2266 -60 -2265
rect -51 -2273 -48 -2250
rect -10 -2231 10 -2228
rect 3923 -2221 3924 -2220
rect 3933 -2228 3936 -2205
rect 3974 -2186 3994 -2183
rect 3974 -2192 3977 -2186
rect 3991 -2192 3994 -2186
rect 3955 -2213 3958 -2210
rect 3955 -2216 3973 -2213
rect 3983 -2223 3986 -2216
rect 3983 -2226 4000 -2223
rect 3905 -2229 3924 -2228
rect 3900 -2231 3924 -2229
rect 3933 -2231 3976 -2228
rect -10 -2237 -7 -2231
rect 7 -2237 10 -2231
rect 3906 -2237 3909 -2231
rect 3997 -2237 4000 -2226
rect -29 -2258 -26 -2255
rect -29 -2261 -11 -2258
rect 3962 -2242 3987 -2239
rect 3997 -2241 4010 -2237
rect 3962 -2244 3965 -2242
rect 3889 -2260 3892 -2257
rect 3897 -2260 3907 -2257
rect 3915 -2257 3918 -2249
rect 3927 -2247 3965 -2244
rect 3997 -2245 4000 -2241
rect 3927 -2257 3930 -2247
rect 3968 -2248 4000 -2245
rect 3968 -2251 3971 -2248
rect 3915 -2260 3930 -2257
rect -1 -2268 2 -2261
rect 3915 -2263 3918 -2260
rect -1 -2271 16 -2268
rect -79 -2274 -60 -2273
rect -84 -2276 -60 -2274
rect -51 -2276 -8 -2273
rect -78 -2282 -75 -2276
rect 13 -2282 16 -2271
rect 3967 -2254 3973 -2251
rect 3906 -2273 3909 -2269
rect 3927 -2270 3932 -2267
rect 3945 -2267 3948 -2263
rect 3992 -2267 3995 -2263
rect 3937 -2270 4001 -2267
rect 3927 -2273 3930 -2270
rect 3900 -2276 3930 -2273
rect 4006 -2281 4010 -2241
rect -22 -2287 3 -2284
rect 13 -2286 26 -2282
rect -22 -2289 -19 -2287
rect -95 -2305 -92 -2302
rect -87 -2305 -77 -2302
rect -69 -2302 -66 -2294
rect -57 -2292 -19 -2289
rect 13 -2290 16 -2286
rect -57 -2302 -54 -2292
rect -16 -2293 16 -2290
rect -16 -2296 -13 -2293
rect -69 -2305 -54 -2302
rect -69 -2308 -66 -2305
rect -17 -2299 -11 -2296
rect -78 -2318 -75 -2314
rect -57 -2315 -52 -2312
rect -39 -2312 -36 -2308
rect 8 -2312 11 -2308
rect -47 -2315 17 -2312
rect -57 -2318 -54 -2315
rect -84 -2321 -54 -2318
rect 22 -2326 26 -2286
rect 401 -2346 424 -2342
rect 405 -2348 424 -2346
rect 401 -2357 405 -2352
rect 420 -2357 424 -2348
rect 437 -2353 461 -2352
rect 437 -2357 453 -2353
rect 457 -2357 461 -2353
rect 437 -2359 461 -2357
rect 443 -2364 447 -2359
rect 412 -2385 416 -2377
rect 412 -2389 424 -2385
rect 420 -2391 424 -2389
rect 451 -2391 455 -2384
rect 395 -2396 413 -2392
rect 420 -2395 444 -2391
rect 451 -2395 461 -2391
rect 395 -2403 402 -2399
rect 420 -2406 424 -2395
rect 451 -2398 455 -2395
rect 443 -2412 447 -2408
rect 437 -2413 462 -2412
rect 437 -2417 457 -2413
rect 437 -2418 462 -2417
rect 401 -2430 405 -2426
rect 401 -2434 417 -2430
rect -86 -2564 -58 -2561
rect -85 -2570 -82 -2564
rect -61 -2565 -58 -2564
rect -61 -2568 10 -2565
rect -102 -2594 -99 -2591
rect -94 -2593 -84 -2590
rect -76 -2590 -73 -2582
rect -46 -2574 -43 -2568
rect -27 -2574 -24 -2568
rect -76 -2593 -55 -2590
rect -76 -2596 -73 -2593
rect -85 -2606 -82 -2602
rect -91 -2608 -67 -2606
rect -91 -2609 -73 -2608
rect -68 -2609 -67 -2608
rect -58 -2616 -55 -2593
rect -17 -2574 3 -2571
rect -17 -2580 -14 -2574
rect 0 -2580 3 -2574
rect -36 -2601 -33 -2598
rect -36 -2604 -18 -2601
rect -8 -2611 -5 -2604
rect 3845 -2606 3873 -2603
rect -8 -2614 9 -2611
rect -86 -2617 -67 -2616
rect -91 -2619 -67 -2617
rect -58 -2619 -15 -2616
rect -85 -2625 -82 -2619
rect 6 -2625 9 -2614
rect 3846 -2612 3849 -2606
rect 3870 -2607 3873 -2606
rect 3870 -2610 3941 -2607
rect -29 -2630 -4 -2627
rect 6 -2629 19 -2625
rect -29 -2632 -26 -2630
rect -102 -2648 -99 -2645
rect -94 -2648 -84 -2645
rect -76 -2645 -73 -2637
rect -64 -2635 -26 -2632
rect 6 -2633 9 -2629
rect -64 -2645 -61 -2635
rect -23 -2636 9 -2633
rect -23 -2639 -20 -2636
rect -76 -2648 -61 -2645
rect -76 -2651 -73 -2648
rect -24 -2642 -18 -2639
rect -85 -2661 -82 -2657
rect -64 -2658 -59 -2655
rect -46 -2655 -43 -2651
rect 1 -2655 4 -2651
rect -54 -2658 10 -2655
rect -64 -2661 -61 -2658
rect -91 -2664 -61 -2661
rect 15 -2669 19 -2629
rect 3829 -2636 3832 -2633
rect 3837 -2635 3847 -2632
rect 3855 -2632 3858 -2624
rect 3885 -2616 3888 -2610
rect 3904 -2616 3907 -2610
rect 3855 -2635 3876 -2632
rect 3855 -2638 3858 -2635
rect 3846 -2648 3849 -2644
rect 3840 -2650 3864 -2648
rect 3840 -2651 3858 -2650
rect 3863 -2651 3864 -2650
rect 3873 -2658 3876 -2635
rect 3914 -2616 3934 -2613
rect 3914 -2622 3917 -2616
rect 3931 -2622 3934 -2616
rect 3895 -2643 3898 -2640
rect 3895 -2646 3913 -2643
rect 3923 -2653 3926 -2646
rect 3923 -2656 3940 -2653
rect 3845 -2659 3864 -2658
rect 3840 -2661 3864 -2659
rect 3873 -2661 3916 -2658
rect 3846 -2667 3849 -2661
rect 3937 -2667 3940 -2656
rect 3902 -2672 3927 -2669
rect 3937 -2671 3950 -2667
rect 3902 -2674 3905 -2672
rect 3829 -2690 3832 -2687
rect 3837 -2690 3847 -2687
rect 3855 -2687 3858 -2679
rect 3867 -2677 3905 -2674
rect 3937 -2675 3940 -2671
rect 3867 -2687 3870 -2677
rect 3908 -2678 3940 -2675
rect 3908 -2681 3911 -2678
rect 3855 -2690 3870 -2687
rect 3855 -2693 3858 -2690
rect 3907 -2684 3913 -2681
rect 3846 -2703 3849 -2699
rect 3867 -2700 3872 -2697
rect 3885 -2697 3888 -2693
rect 3932 -2697 3935 -2693
rect 3877 -2700 3941 -2697
rect 3867 -2703 3870 -2700
rect 3840 -2706 3870 -2703
rect 389 -2712 412 -2708
rect 3946 -2711 3950 -2671
rect 393 -2714 412 -2712
rect 389 -2723 393 -2718
rect 408 -2723 412 -2714
rect 425 -2719 449 -2718
rect 425 -2723 441 -2719
rect 445 -2723 449 -2719
rect 425 -2725 449 -2723
rect 431 -2730 435 -2725
rect 400 -2751 404 -2743
rect 400 -2755 412 -2751
rect 408 -2757 412 -2755
rect 439 -2757 443 -2750
rect 383 -2762 401 -2758
rect 408 -2761 432 -2757
rect 439 -2761 449 -2757
rect 383 -2769 390 -2765
rect 408 -2772 412 -2761
rect 439 -2764 443 -2761
rect 431 -2778 435 -2774
rect 425 -2779 450 -2778
rect 425 -2783 445 -2779
rect 425 -2784 450 -2783
rect 389 -2796 393 -2792
rect 389 -2800 405 -2796
rect 3802 -3142 3830 -3139
rect 3803 -3148 3806 -3142
rect 3827 -3143 3830 -3142
rect 3827 -3146 3898 -3143
rect 3786 -3172 3789 -3169
rect 3794 -3171 3804 -3168
rect 3812 -3168 3815 -3160
rect 3842 -3152 3845 -3146
rect 3861 -3152 3864 -3146
rect 3812 -3171 3833 -3168
rect 3812 -3174 3815 -3171
rect 3803 -3184 3806 -3180
rect 3797 -3186 3821 -3184
rect 3797 -3187 3815 -3186
rect 3820 -3187 3821 -3186
rect 3830 -3194 3833 -3171
rect 3871 -3152 3891 -3149
rect 3871 -3158 3874 -3152
rect 3888 -3158 3891 -3152
rect 3852 -3179 3855 -3176
rect 3852 -3182 3870 -3179
rect 3880 -3189 3883 -3182
rect 3880 -3192 3897 -3189
rect 3802 -3195 3821 -3194
rect 3797 -3197 3821 -3195
rect 3830 -3197 3873 -3194
rect 3803 -3203 3806 -3197
rect 3894 -3203 3897 -3192
rect 3859 -3208 3884 -3205
rect 3894 -3207 3907 -3203
rect 3859 -3210 3862 -3208
rect 3786 -3226 3789 -3223
rect 3794 -3226 3804 -3223
rect 3812 -3223 3815 -3215
rect 3824 -3213 3862 -3210
rect 3894 -3211 3897 -3207
rect 3824 -3223 3827 -3213
rect 3865 -3214 3897 -3211
rect 3865 -3217 3868 -3214
rect 3812 -3226 3827 -3223
rect 3812 -3229 3815 -3226
rect 3864 -3220 3870 -3217
rect 3803 -3239 3806 -3235
rect 3824 -3236 3829 -3233
rect 3842 -3233 3845 -3229
rect 3889 -3233 3892 -3229
rect 3834 -3236 3898 -3233
rect 3824 -3239 3827 -3236
rect 3797 -3242 3827 -3239
rect 3903 -3247 3907 -3207
<< m2contact >>
rect 3852 -1397 3857 -1392
rect 3852 -1451 3857 -1446
rect -110 -1534 -105 -1529
rect -110 -1588 -105 -1583
rect -119 -1893 -114 -1888
rect -119 -1947 -114 -1942
rect 3892 -2207 3897 -2202
rect -92 -2252 -87 -2247
rect 3892 -2261 3897 -2256
rect -92 -2306 -87 -2301
rect -99 -2595 -94 -2590
rect -99 -2649 -94 -2644
rect 3832 -2637 3837 -2632
rect 3832 -2691 3837 -2686
rect 3789 -3173 3794 -3168
rect 3789 -3227 3794 -3222
<< pm12contact >>
rect 3908 -1414 3913 -1409
rect 3917 -1415 3922 -1410
rect -54 -1551 -49 -1546
rect -45 -1552 -40 -1547
rect 1601 -1680 1607 -1674
rect 1651 -1679 1657 -1673
rect 1701 -1679 1707 -1673
rect 1748 -1679 1754 -1673
rect -63 -1910 -58 -1905
rect -54 -1911 -49 -1906
rect 2071 -1893 2076 -1888
rect 2109 -1893 2114 -1888
rect 2153 -1893 2158 -1888
rect 2191 -1893 2196 -1888
rect 2237 -1891 2242 -1886
rect 1538 -1955 1543 -1950
rect 1566 -1955 1571 -1950
rect 1593 -1955 1598 -1950
rect 1632 -1955 1637 -1950
rect 1660 -1955 1665 -1950
rect 1687 -1955 1692 -1950
rect 1727 -1954 1732 -1949
rect 1755 -1954 1760 -1949
rect 1782 -1954 1787 -1949
rect 1818 -1954 1823 -1949
rect 3948 -2224 3953 -2219
rect 3957 -2225 3962 -2220
rect -36 -2269 -31 -2264
rect -27 -2270 -22 -2265
rect -43 -2612 -38 -2607
rect -34 -2613 -29 -2608
rect 3888 -2654 3893 -2649
rect 3897 -2655 3902 -2650
rect 3845 -3190 3850 -3185
rect 3854 -3191 3859 -3186
<< metal2 >>
rect 3853 -1403 3856 -1397
rect 3853 -1406 3890 -1403
rect 3887 -1409 3890 -1406
rect 3887 -1412 3908 -1409
rect 3917 -1425 3920 -1415
rect 3854 -1428 3920 -1425
rect 3854 -1446 3857 -1428
rect -109 -1540 -106 -1534
rect -109 -1543 -72 -1540
rect -75 -1546 -72 -1543
rect -75 -1549 -54 -1546
rect -45 -1562 -42 -1552
rect -108 -1565 -42 -1562
rect -108 -1583 -105 -1565
rect 1591 -1680 1601 -1674
rect 1641 -1679 1651 -1673
rect 1691 -1679 1701 -1673
rect 1738 -1679 1748 -1673
rect 2068 -1893 2071 -1888
rect 2106 -1893 2109 -1888
rect 2150 -1893 2153 -1888
rect 2188 -1893 2191 -1888
rect 2234 -1891 2237 -1886
rect -118 -1899 -115 -1893
rect -118 -1902 -81 -1899
rect -84 -1905 -81 -1902
rect -84 -1908 -63 -1905
rect -54 -1921 -51 -1911
rect -117 -1924 -51 -1921
rect -117 -1942 -114 -1924
rect 1534 -1955 1538 -1950
rect 1562 -1955 1566 -1950
rect 1589 -1955 1593 -1950
rect 1628 -1955 1632 -1950
rect 1656 -1955 1660 -1950
rect 1683 -1955 1687 -1950
rect 1723 -1954 1727 -1949
rect 1751 -1954 1755 -1949
rect 1778 -1954 1782 -1949
rect 1814 -1954 1818 -1949
rect 3893 -2213 3896 -2207
rect 3893 -2216 3930 -2213
rect 3927 -2219 3930 -2216
rect 3927 -2222 3948 -2219
rect 3957 -2235 3960 -2225
rect 3894 -2238 3960 -2235
rect -91 -2258 -88 -2252
rect 3894 -2256 3897 -2238
rect -91 -2261 -54 -2258
rect -57 -2264 -54 -2261
rect -57 -2267 -36 -2264
rect -27 -2280 -24 -2270
rect -90 -2283 -24 -2280
rect -90 -2301 -87 -2283
rect -98 -2601 -95 -2595
rect -98 -2604 -61 -2601
rect -64 -2607 -61 -2604
rect -64 -2610 -43 -2607
rect -34 -2623 -31 -2613
rect -97 -2626 -31 -2623
rect -97 -2644 -94 -2626
rect 3833 -2643 3836 -2637
rect 3833 -2646 3870 -2643
rect 3867 -2649 3870 -2646
rect 3867 -2652 3888 -2649
rect 3897 -2665 3900 -2655
rect 3834 -2668 3900 -2665
rect 3834 -2686 3837 -2668
rect 3790 -3179 3793 -3173
rect 3790 -3182 3827 -3179
rect 3824 -3185 3827 -3182
rect 3824 -3188 3845 -3185
rect 3854 -3201 3857 -3191
rect 3791 -3204 3857 -3201
rect 3791 -3222 3794 -3204
<< m123contact >>
rect 3860 -1366 3865 -1361
rect 3860 -1419 3865 -1414
rect 3878 -1415 3883 -1410
rect 3892 -1460 3897 -1455
rect -102 -1503 -97 -1498
rect -102 -1556 -97 -1551
rect -84 -1552 -79 -1547
rect -70 -1597 -65 -1592
rect -111 -1862 -106 -1857
rect -111 -1915 -106 -1910
rect -93 -1911 -88 -1906
rect -79 -1956 -74 -1951
rect 3900 -2176 3905 -2171
rect -84 -2221 -79 -2216
rect 3900 -2229 3905 -2224
rect 3918 -2225 3923 -2220
rect -84 -2274 -79 -2269
rect -66 -2270 -61 -2265
rect 3932 -2270 3937 -2265
rect -52 -2315 -47 -2310
rect -91 -2564 -86 -2559
rect 3840 -2606 3845 -2601
rect -91 -2617 -86 -2612
rect -73 -2613 -68 -2608
rect -59 -2658 -54 -2653
rect 3840 -2659 3845 -2654
rect 3858 -2655 3863 -2650
rect 3872 -2700 3877 -2695
rect 3797 -3142 3802 -3137
rect 3797 -3195 3802 -3190
rect 3815 -3191 3820 -3186
rect 3829 -3236 3834 -3231
<< metal3 >>
rect 3860 -1414 3863 -1366
rect 3883 -1415 3895 -1412
rect 3892 -1455 3895 -1415
rect -102 -1551 -99 -1503
rect -79 -1552 -67 -1549
rect -70 -1592 -67 -1552
rect -111 -1910 -108 -1862
rect -88 -1911 -76 -1908
rect -79 -1951 -76 -1911
rect -84 -2269 -81 -2221
rect 3900 -2224 3903 -2176
rect 3923 -2225 3935 -2222
rect 3932 -2265 3935 -2225
rect -61 -2270 -49 -2267
rect -52 -2310 -49 -2270
rect -91 -2612 -88 -2564
rect -68 -2613 -56 -2610
rect -59 -2653 -56 -2613
rect 3840 -2654 3843 -2606
rect 3863 -2655 3875 -2652
rect 3872 -2695 3875 -2655
rect 3797 -3190 3800 -3142
rect 3820 -3191 3832 -3188
rect 3829 -3231 3832 -3191
<< labels >>
rlabel metal1 1538 -1839 1542 -1835 1 pdr1
rlabel metal2 1534 -1955 1538 -1950 2 prop_1
rlabel metal1 1546 -1949 1550 -1944 1 prop1_car0
rlabel metal1 1566 -1840 1570 -1835 1 prop1_car0
rlabel metal2 1562 -1955 1566 -1950 1 carry_0
rlabel metal1 1574 -1949 1578 -1944 1 clock_car0
rlabel metal1 1593 -1840 1597 -1835 1 clock_car0
rlabel metal2 1589 -1955 1593 -1950 1 clock_in
rlabel metal1 1601 -1949 1605 -1944 1 gnd!
rlabel metal1 1632 -1840 1636 -1835 1 pdr2
rlabel metal2 1628 -1955 1632 -1950 1 prop_2
rlabel metal1 1640 -1949 1644 -1944 1 pdr1
rlabel metal1 1660 -1840 1664 -1835 1 pdr1
rlabel metal2 1656 -1955 1660 -1950 1 gen_1
rlabel metal1 1668 -1949 1672 -1944 1 clock_car0
rlabel metal1 1687 -1840 1691 -1835 1 pdr3
rlabel metal2 1683 -1955 1687 -1950 1 prop_3
rlabel metal1 1695 -1949 1699 -1944 1 pdr2
rlabel metal1 1727 -1839 1731 -1834 1 pdr2
rlabel metal2 1723 -1954 1727 -1949 1 gen_2
rlabel metal1 1735 -1948 1739 -1943 1 clock_car0
rlabel metal1 1755 -1839 1759 -1834 1 pdr4
rlabel metal2 1751 -1954 1755 -1949 1 prop_4
rlabel metal1 1763 -1948 1767 -1943 1 pdr3
rlabel metal1 1782 -1839 1786 -1834 1 pdr3
rlabel metal2 1778 -1954 1782 -1949 1 gen_3
rlabel metal1 1790 -1948 1794 -1943 1 clock_car0
rlabel metal1 1818 -1839 1822 -1834 1 pdr4
rlabel metal2 1814 -1954 1818 -1949 1 gen_4
rlabel metal1 1826 -1948 1830 -1943 7 clock_car0
rlabel metal1 1602 -1592 1606 -1587 5 vdd!
rlabel metal1 1652 -1591 1656 -1586 5 vdd!
rlabel metal1 1702 -1591 1706 -1586 5 vdd!
rlabel metal1 1749 -1591 1753 -1586 5 vdd!
rlabel metal2 1591 -1680 1597 -1674 2 clock_in
rlabel metal2 1641 -1679 1647 -1673 1 clock_in
rlabel metal2 1691 -1679 1697 -1673 1 clock_in
rlabel metal2 1738 -1679 1743 -1673 1 clock_in
rlabel metal1 1610 -1671 1614 -1666 1 pdr1
rlabel metal1 1660 -1670 1664 -1666 1 pdr2
rlabel metal1 1710 -1670 1714 -1666 1 pdr3
rlabel metal1 1757 -1670 1761 -1666 1 pdr4
rlabel metal1 2196 -1929 2200 -1925 1 gnd!
rlabel metal1 2192 -1825 2197 -1821 5 vdd!
rlabel metal2 2068 -1893 2071 -1888 1 pdr1
rlabel metal2 2106 -1893 2109 -1888 1 pdr2
rlabel metal2 2150 -1893 2153 -1888 1 pdr3
rlabel metal2 2188 -1893 2191 -1888 1 pdr4
rlabel metal1 2079 -1893 2083 -1888 1 c1
rlabel metal1 2117 -1893 2121 -1888 1 c2
rlabel metal1 2161 -1893 2165 -1888 1 c3
rlabel metal1 2199 -1893 2203 -1888 1 c4
rlabel metal1 2242 -1927 2246 -1923 1 gnd!
rlabel metal1 2238 -1823 2243 -1819 5 vdd!
rlabel metal2 2234 -1891 2237 -1886 1 clk_org
rlabel metal1 2245 -1891 2249 -1886 1 clock_in
rlabel metal1 2071 -1825 2075 -1821 5 vdd!
rlabel metal1 2109 -1825 2113 -1821 5 vdd!
rlabel metal1 2153 -1825 2157 -1821 5 vdd!
rlabel metal1 2157 -1929 2161 -1925 1 gnd!
rlabel metal1 2120 -1929 2124 -1925 1 gnd!
rlabel metal1 2080 -1929 2084 -1925 1 gnd!
rlabel metal1 401 -1703 401 -1703 5 vdd
rlabel metal1 402 -1790 402 -1790 1 gnd
rlabel metal1 434 -1772 434 -1772 1 gnd
rlabel metal1 431 -1715 431 -1715 5 vdd
rlabel metal1 403 -2053 403 -2053 5 vdd
rlabel metal1 404 -2140 404 -2140 1 gnd
rlabel metal1 436 -2122 436 -2122 1 gnd
rlabel metal1 433 -2065 433 -2065 5 vdd
rlabel metal1 411 -2345 411 -2345 5 vdd
rlabel metal1 412 -2432 412 -2432 1 gnd
rlabel metal1 444 -2414 444 -2414 1 gnd
rlabel metal1 441 -2357 441 -2357 5 vdd
rlabel metal1 399 -2711 399 -2711 5 vdd
rlabel metal1 400 -2798 400 -2798 1 gnd
rlabel metal1 432 -2780 432 -2780 1 gnd
rlabel metal1 429 -2723 429 -2723 5 vdd
rlabel metal1 386 -1752 386 -1752 3 q_a1
rlabel metal1 388 -1759 388 -1759 3 q_b1
rlabel metal1 450 -1752 450 -1752 1 gen_1
rlabel metal1 389 -2103 389 -2103 1 q_a2
rlabel metal1 389 -2110 389 -2110 1 q_b2
rlabel metal1 452 -2101 452 -2101 1 gen_2
rlabel metal1 396 -2395 396 -2395 1 q_b3
rlabel metal1 398 -2402 398 -2402 1 q_a3
rlabel metal1 459 -2393 459 -2393 1 gen_3
rlabel metal1 384 -2760 384 -2760 3 q_a4
rlabel metal1 384 -2766 384 -2766 3 q_b4
rlabel metal1 447 -2759 447 -2759 1 gen_4
rlabel metal1 -84 -1603 -80 -1600 1 gnd
rlabel metal1 -34 -1597 -31 -1595 1 gnd
rlabel metal1 -86 -1547 -85 -1545 1 gnd
rlabel metal1 -90 -1503 -87 -1501 5 vdd
rlabel metal1 -89 -1557 -86 -1555 1 vdd
rlabel metal1 -93 -1962 -89 -1959 1 gnd
rlabel metal1 -43 -1956 -40 -1954 1 gnd
rlabel metal1 -95 -1906 -94 -1904 1 gnd
rlabel metal1 -99 -1862 -96 -1860 5 vdd
rlabel metal1 -98 -1916 -95 -1914 1 vdd
rlabel metal1 -66 -2321 -62 -2318 1 gnd
rlabel metal1 -16 -2315 -13 -2313 1 gnd
rlabel metal1 -68 -2265 -67 -2263 1 gnd
rlabel metal1 -72 -2221 -69 -2219 5 vdd
rlabel metal1 -71 -2275 -68 -2273 1 vdd
rlabel metal1 -73 -2664 -69 -2661 1 gnd
rlabel metal1 -23 -2658 -20 -2656 1 gnd
rlabel metal1 -75 -2608 -74 -2606 1 gnd
rlabel metal1 -79 -2564 -76 -2562 5 vdd
rlabel metal1 -78 -2618 -75 -2616 1 vdd
rlabel metal1 3878 -1466 3882 -1463 1 gnd
rlabel metal1 3928 -1460 3931 -1458 1 gnd
rlabel metal1 3876 -1410 3877 -1408 1 gnd
rlabel metal1 3872 -1366 3875 -1364 5 vdd
rlabel metal1 3873 -1420 3876 -1418 1 vdd
rlabel metal1 3918 -2276 3922 -2273 1 gnd
rlabel metal1 3968 -2270 3971 -2268 1 gnd
rlabel metal1 3916 -2220 3917 -2218 1 gnd
rlabel metal1 3912 -2176 3915 -2174 5 vdd
rlabel metal1 3913 -2230 3916 -2228 1 vdd
rlabel metal1 3858 -2706 3862 -2703 1 gnd
rlabel metal1 3908 -2700 3911 -2698 1 gnd
rlabel metal1 3856 -2650 3857 -2648 1 gnd
rlabel metal1 3852 -2606 3855 -2604 5 vdd
rlabel metal1 3853 -2660 3856 -2658 1 vdd
rlabel metal1 -112 -1531 -112 -1531 1 q_a1
rlabel metal1 -112 -1585 -112 -1585 1 q_b1
rlabel metal1 4 -1566 4 -1566 1 prop_1
rlabel metal1 -121 -1890 -121 -1890 3 q_a2
rlabel metal1 -121 -1945 -121 -1945 3 q_b2
rlabel metal1 -3 -1924 -3 -1924 1 prop_2
rlabel metal1 -93 -2249 -93 -2249 1 q_a3
rlabel metal1 -93 -2303 -93 -2303 1 q_b3
rlabel metal1 24 -2284 24 -2284 1 prop_3
rlabel metal1 -101 -2593 -101 -2593 1 q_a4
rlabel metal1 -101 -2646 -101 -2646 1 q_b4
rlabel metal1 18 -2627 18 -2627 1 prop_4
rlabel metal1 3850 -1394 3850 -1394 1 carry_0
rlabel metal1 3850 -1448 3850 -1448 1 prop_1
rlabel metal1 3969 -1429 3969 -1429 1 s1
rlabel metal1 3891 -2205 3891 -2205 1 c1
rlabel metal1 3890 -2259 3890 -2259 1 prop_2
rlabel metal1 4009 -2240 4009 -2240 7 s2
rlabel metal1 3830 -2634 3830 -2634 1 c2
rlabel metal1 3830 -2689 3830 -2689 1 prop_3
rlabel metal1 3949 -2669 3949 -2669 1 s3
rlabel metal1 3815 -3242 3819 -3239 1 gnd
rlabel metal1 3865 -3236 3868 -3234 1 gnd
rlabel metal1 3813 -3186 3814 -3184 1 gnd
rlabel metal1 3809 -3142 3812 -3140 5 vdd
rlabel metal1 3810 -3196 3813 -3194 1 vdd
rlabel metal1 3905 -3205 3905 -3205 1 s4
rlabel metal1 3787 -3224 3787 -3224 1 prop_4
rlabel metal1 3787 -3171 3787 -3171 1 c3
<< end >>
