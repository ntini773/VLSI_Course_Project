magic
tech scmos
timestamp 1732004421
<< nwell >>
rect 112 -313 136 -251
rect 162 -312 186 -250
rect 212 -312 236 -250
rect 259 -312 283 -250
rect 581 -534 605 -482
rect 619 -534 643 -482
rect 663 -534 687 -482
rect 701 -534 725 -482
rect 747 -532 771 -480
<< ntransistor >>
rect 59 -593 61 -493
rect 87 -593 89 -493
rect 114 -593 116 -493
rect 153 -593 155 -493
rect 181 -593 183 -493
rect 208 -593 210 -493
rect 248 -592 250 -492
rect 276 -592 278 -492
rect 303 -592 305 -492
rect 339 -592 341 -492
rect 592 -566 594 -546
rect 630 -566 632 -546
rect 674 -566 676 -546
rect 712 -566 714 -546
rect 758 -564 760 -544
<< ptransistor >>
rect 123 -307 125 -257
rect 173 -306 175 -256
rect 223 -306 225 -256
rect 270 -306 272 -256
rect 592 -528 594 -488
rect 630 -528 632 -488
rect 674 -528 676 -488
rect 712 -528 714 -488
rect 758 -526 760 -486
<< ndiffusion >>
rect 58 -593 59 -493
rect 61 -593 62 -493
rect 86 -593 87 -493
rect 89 -593 90 -493
rect 113 -593 114 -493
rect 116 -593 117 -493
rect 152 -593 153 -493
rect 155 -593 156 -493
rect 180 -593 181 -493
rect 183 -593 184 -493
rect 207 -593 208 -493
rect 210 -593 211 -493
rect 247 -592 248 -492
rect 250 -592 251 -492
rect 275 -592 276 -492
rect 278 -592 279 -492
rect 302 -592 303 -492
rect 305 -592 306 -492
rect 338 -592 339 -492
rect 341 -592 342 -492
rect 591 -566 592 -546
rect 594 -566 595 -546
rect 629 -566 630 -546
rect 632 -566 633 -546
rect 673 -566 674 -546
rect 676 -566 677 -546
rect 711 -566 712 -546
rect 714 -566 715 -546
rect 757 -564 758 -544
rect 760 -564 761 -544
<< pdiffusion >>
rect 122 -307 123 -257
rect 125 -307 126 -257
rect 172 -306 173 -256
rect 175 -306 176 -256
rect 222 -306 223 -256
rect 225 -306 226 -256
rect 269 -306 270 -256
rect 272 -306 273 -256
rect 591 -528 592 -488
rect 594 -528 595 -488
rect 629 -528 630 -488
rect 632 -528 633 -488
rect 673 -528 674 -488
rect 676 -528 677 -488
rect 711 -528 712 -488
rect 714 -528 715 -488
rect 757 -526 758 -486
rect 760 -526 761 -486
<< ndcontact >>
rect 54 -593 58 -493
rect 62 -593 66 -493
rect 82 -593 86 -493
rect 90 -593 94 -493
rect 109 -593 113 -493
rect 117 -593 121 -493
rect 148 -593 152 -493
rect 156 -593 160 -493
rect 176 -593 180 -493
rect 184 -593 188 -493
rect 203 -593 207 -493
rect 211 -593 215 -493
rect 243 -592 247 -492
rect 251 -592 255 -492
rect 271 -592 275 -492
rect 279 -592 283 -492
rect 298 -592 302 -492
rect 306 -592 310 -492
rect 334 -592 338 -492
rect 342 -592 346 -492
rect 587 -566 591 -546
rect 595 -566 599 -546
rect 625 -566 629 -546
rect 633 -566 637 -546
rect 669 -566 673 -546
rect 677 -566 681 -546
rect 707 -566 711 -546
rect 715 -566 719 -546
rect 753 -564 757 -544
rect 761 -564 765 -544
<< pdcontact >>
rect 118 -307 122 -257
rect 126 -307 130 -257
rect 168 -306 172 -256
rect 176 -306 180 -256
rect 218 -306 222 -256
rect 226 -306 230 -256
rect 265 -306 269 -256
rect 273 -306 277 -256
rect 587 -528 591 -488
rect 595 -528 599 -488
rect 625 -528 629 -488
rect 633 -528 637 -488
rect 669 -528 673 -488
rect 677 -528 681 -488
rect 707 -528 711 -488
rect 715 -528 719 -488
rect 753 -526 757 -486
rect 761 -526 765 -486
<< nsubstratencontact >>
rect 113 -251 117 -246
rect 163 -250 167 -245
rect 213 -250 217 -245
rect 260 -250 264 -245
rect 582 -482 586 -478
rect 620 -482 624 -478
rect 664 -482 668 -478
rect 702 -482 706 -478
rect 748 -480 752 -476
<< polysilicon >>
rect 123 -257 125 -254
rect 173 -256 175 -253
rect 223 -256 225 -253
rect 270 -256 272 -253
rect 123 -330 125 -307
rect 173 -329 175 -306
rect 223 -329 225 -306
rect 270 -329 272 -306
rect 592 -488 594 -485
rect 630 -488 632 -485
rect 674 -488 676 -485
rect 712 -488 714 -485
rect 758 -486 760 -483
rect 59 -493 61 -490
rect 87 -493 89 -490
rect 114 -493 116 -490
rect 153 -493 155 -490
rect 181 -493 183 -490
rect 208 -493 210 -490
rect 248 -492 250 -489
rect 276 -492 278 -489
rect 303 -492 305 -489
rect 339 -492 341 -489
rect 592 -546 594 -528
rect 630 -546 632 -528
rect 674 -546 676 -528
rect 712 -546 714 -528
rect 758 -544 760 -526
rect 592 -570 594 -566
rect 630 -570 632 -566
rect 674 -570 676 -566
rect 712 -570 714 -566
rect 758 -568 760 -564
rect 59 -605 61 -593
rect 87 -605 89 -593
rect 114 -605 116 -593
rect 153 -605 155 -593
rect 181 -605 183 -593
rect 208 -605 210 -593
rect 248 -604 250 -592
rect 276 -604 278 -592
rect 303 -604 305 -592
rect 339 -604 341 -592
<< metal1 >>
rect 118 -246 122 -237
rect 168 -245 172 -236
rect 218 -245 222 -236
rect 265 -245 269 -236
rect 112 -251 113 -246
rect 117 -251 136 -246
rect 162 -250 163 -245
rect 167 -250 186 -245
rect 212 -250 213 -245
rect 217 -250 236 -245
rect 259 -250 260 -245
rect 264 -250 283 -245
rect 118 -257 122 -251
rect 168 -256 172 -250
rect 218 -256 222 -250
rect 265 -256 269 -250
rect 126 -321 130 -307
rect 176 -320 180 -306
rect 226 -320 230 -306
rect 273 -320 277 -306
rect 587 -475 607 -471
rect 618 -475 649 -471
rect 661 -475 689 -471
rect 699 -475 720 -471
rect 736 -473 766 -469
rect 587 -478 591 -475
rect 625 -478 629 -475
rect 669 -478 673 -475
rect 707 -478 711 -475
rect 753 -476 757 -473
rect 581 -482 582 -478
rect 586 -482 591 -478
rect 619 -482 620 -478
rect 624 -482 629 -478
rect 663 -482 664 -478
rect 668 -482 673 -478
rect 701 -482 702 -478
rect 706 -482 711 -478
rect 747 -480 748 -476
rect 752 -480 757 -476
rect 54 -493 58 -485
rect 82 -493 86 -485
rect 109 -493 113 -485
rect 148 -493 152 -485
rect 176 -493 180 -485
rect 203 -493 207 -485
rect 243 -492 247 -484
rect 271 -492 275 -484
rect 298 -492 302 -484
rect 334 -492 338 -484
rect 587 -488 591 -482
rect 625 -488 629 -482
rect 669 -488 673 -482
rect 707 -488 711 -482
rect 753 -486 757 -480
rect 595 -546 599 -528
rect 633 -546 637 -528
rect 677 -546 681 -528
rect 715 -546 719 -528
rect 761 -544 765 -526
rect 587 -575 591 -566
rect 625 -575 629 -566
rect 669 -575 673 -566
rect 707 -575 711 -566
rect 753 -573 757 -564
rect 587 -579 607 -575
rect 618 -579 649 -575
rect 661 -579 689 -575
rect 699 -579 716 -575
rect 736 -577 762 -573
rect 62 -599 66 -593
rect 90 -599 94 -593
rect 117 -599 121 -593
rect 156 -599 160 -593
rect 184 -599 188 -593
rect 211 -599 215 -593
rect 251 -598 255 -592
rect 279 -598 283 -592
rect 306 -598 310 -592
rect 342 -598 346 -592
<< pm12contact >>
rect 117 -330 123 -324
rect 167 -329 173 -323
rect 217 -329 223 -323
rect 264 -329 270 -323
rect 587 -543 592 -538
rect 625 -543 630 -538
rect 669 -543 674 -538
rect 707 -543 712 -538
rect 753 -541 758 -536
rect 54 -605 59 -600
rect 82 -605 87 -600
rect 109 -605 114 -600
rect 148 -605 153 -600
rect 176 -605 181 -600
rect 203 -605 208 -600
rect 243 -604 248 -599
rect 271 -604 276 -599
rect 298 -604 303 -599
rect 334 -604 339 -599
<< metal2 >>
rect 107 -330 117 -324
rect 157 -329 167 -323
rect 207 -329 217 -323
rect 254 -329 264 -323
rect 584 -543 587 -538
rect 622 -543 625 -538
rect 666 -543 669 -538
rect 704 -543 707 -538
rect 750 -541 753 -536
rect 50 -605 54 -600
rect 78 -605 82 -600
rect 105 -605 109 -600
rect 144 -605 148 -600
rect 172 -605 176 -600
rect 199 -605 203 -600
rect 239 -604 243 -599
rect 267 -604 271 -599
rect 294 -604 298 -599
rect 330 -604 334 -599
<< labels >>
rlabel metal1 54 -489 58 -485 1 pdr1
rlabel metal2 50 -605 54 -600 2 prop_1
rlabel metal1 62 -599 66 -594 1 prop1_car0
rlabel metal1 82 -490 86 -485 1 prop1_car0
rlabel metal2 78 -605 82 -600 1 carry_0
rlabel metal1 90 -599 94 -594 1 clock_car0
rlabel metal1 109 -490 113 -485 1 clock_car0
rlabel metal2 105 -605 109 -600 1 clock_in
rlabel metal1 117 -599 121 -594 1 gnd!
rlabel metal1 148 -490 152 -485 1 pdr2
rlabel metal2 144 -605 148 -600 1 prop_2
rlabel metal1 156 -599 160 -594 1 pdr1
rlabel metal1 176 -490 180 -485 1 pdr1
rlabel metal2 172 -605 176 -600 1 gen_1
rlabel metal1 184 -599 188 -594 1 clock_car0
rlabel metal1 203 -490 207 -485 1 pdr3
rlabel metal2 199 -605 203 -600 1 prop_3
rlabel metal1 211 -599 215 -594 1 pdr2
rlabel metal1 243 -489 247 -484 1 pdr2
rlabel metal2 239 -604 243 -599 1 gen_2
rlabel metal1 251 -598 255 -593 1 clock_car0
rlabel metal1 271 -489 275 -484 1 pdr4
rlabel metal2 267 -604 271 -599 1 prop_4
rlabel metal1 279 -598 283 -593 1 pdr3
rlabel metal1 298 -489 302 -484 1 pdr3
rlabel metal2 294 -604 298 -599 1 gen_3
rlabel metal1 306 -598 310 -593 1 clock_car0
rlabel metal1 334 -489 338 -484 1 pdr4
rlabel metal2 330 -604 334 -599 1 gen_4
rlabel metal1 342 -598 346 -593 7 clock_car0
rlabel metal1 118 -242 122 -237 5 vdd!
rlabel metal1 168 -241 172 -236 5 vdd!
rlabel metal1 218 -241 222 -236 5 vdd!
rlabel metal1 265 -241 269 -236 5 vdd!
rlabel metal2 107 -330 113 -324 2 clock_in
rlabel metal2 157 -329 163 -323 1 clock_in
rlabel metal2 207 -329 213 -323 1 clock_in
rlabel metal2 254 -329 259 -323 1 clock_in
rlabel metal1 126 -321 130 -316 1 pdr1
rlabel metal1 176 -320 180 -316 1 pdr2
rlabel metal1 226 -320 230 -316 1 pdr3
rlabel metal1 273 -320 277 -316 1 pdr4
rlabel metal1 712 -579 716 -575 1 gnd!
rlabel metal1 708 -475 713 -471 5 vdd!
rlabel metal2 584 -543 587 -538 1 pdr1
rlabel metal2 622 -543 625 -538 1 pdr2
rlabel metal2 666 -543 669 -538 1 pdr3
rlabel metal2 704 -543 707 -538 1 pdr4
rlabel metal1 595 -543 599 -538 1 c1
rlabel metal1 633 -543 637 -538 1 c2
rlabel metal1 677 -543 681 -538 1 c3
rlabel metal1 715 -543 719 -538 1 c4
rlabel metal1 758 -577 762 -573 1 gnd!
rlabel metal1 754 -473 759 -469 5 vdd!
rlabel metal2 750 -541 753 -536 1 clk_org
rlabel metal1 761 -541 765 -536 1 clock_in
rlabel metal1 587 -475 591 -471 5 vdd!
rlabel metal1 625 -475 629 -471 5 vdd!
rlabel metal1 669 -475 673 -471 5 vdd!
rlabel metal1 673 -579 677 -575 1 gnd!
rlabel metal1 636 -579 640 -575 1 gnd!
rlabel metal1 596 -579 600 -575 1 gnd!
<< end >>
