magic
tech scmos
timestamp 1732057892
<< nwell >>
rect 2070 -698 2094 -674
rect 2109 -684 2143 -678
rect 2109 -714 2171 -684
rect 2137 -720 2171 -714
rect 2070 -753 2094 -729
rect 2210 -745 2242 -708
rect 2248 -745 2274 -708
rect 2292 -745 2318 -708
rect 2337 -745 2363 -708
rect 2386 -745 2410 -713
rect 2224 -849 2256 -812
rect 2262 -849 2288 -812
rect 2306 -849 2332 -812
rect 2351 -849 2377 -812
rect 2391 -849 2415 -817
rect 957 -916 994 -884
rect 1064 -916 1101 -884
rect 1166 -916 1203 -884
rect 1263 -916 1300 -884
rect 1367 -915 1404 -883
rect 1469 -915 1506 -883
rect 1565 -915 1602 -883
rect 1664 -915 1701 -883
rect 957 -948 994 -922
rect 1064 -948 1101 -922
rect 1166 -948 1203 -922
rect 1263 -948 1300 -922
rect 1367 -947 1404 -921
rect 1469 -947 1506 -921
rect 1565 -947 1602 -921
rect 1664 -947 1701 -921
rect 957 -992 994 -966
rect 1064 -992 1101 -966
rect 1166 -992 1203 -966
rect 1263 -992 1300 -966
rect 1367 -991 1404 -965
rect 1469 -991 1506 -965
rect 1565 -991 1602 -965
rect 1664 -991 1701 -965
rect 2087 -968 2123 -940
rect 2081 -974 2123 -968
rect 2081 -1002 2117 -974
rect 2377 -978 2409 -941
rect 2415 -978 2441 -941
rect 2459 -978 2485 -941
rect 2504 -978 2530 -941
rect 2552 -978 2576 -946
rect 957 -1037 994 -1011
rect 1064 -1037 1101 -1011
rect 1166 -1037 1203 -1011
rect 1263 -1037 1300 -1011
rect 1367 -1036 1404 -1010
rect 1469 -1036 1506 -1010
rect 1565 -1036 1602 -1010
rect 1664 -1036 1701 -1010
rect 2256 -1016 2292 -988
rect 2077 -1041 2101 -1017
rect 2132 -1041 2156 -1017
rect 2250 -1022 2292 -1016
rect 2250 -1050 2286 -1022
rect 1705 -1093 1729 -1069
rect 1744 -1079 1778 -1073
rect 1744 -1109 1806 -1079
rect 2246 -1089 2270 -1065
rect 2301 -1089 2325 -1065
rect 1772 -1115 1806 -1109
rect 1705 -1148 1729 -1124
rect 2571 -1136 2603 -1099
rect 2609 -1136 2635 -1099
rect 2653 -1136 2679 -1099
rect 2698 -1136 2724 -1099
rect 2745 -1136 2769 -1104
rect 2439 -1174 2475 -1146
rect 2433 -1180 2475 -1174
rect 1706 -1225 1730 -1201
rect 1745 -1211 1779 -1205
rect 2433 -1208 2469 -1180
rect 1745 -1241 1807 -1211
rect 1773 -1247 1807 -1241
rect 1706 -1280 1730 -1256
rect 2050 -1263 2102 -1239
rect 2429 -1247 2453 -1223
rect 2484 -1247 2508 -1223
rect 2217 -1306 2269 -1282
rect 2399 -1313 2451 -1289
rect 1709 -1369 1733 -1345
rect 1748 -1355 1782 -1349
rect 1748 -1385 1810 -1355
rect 1776 -1391 1810 -1385
rect 1709 -1424 1733 -1400
rect 2685 -1437 2709 -1385
rect 2732 -1441 2764 -1404
rect 2770 -1441 2796 -1404
rect 2814 -1441 2840 -1404
rect 2859 -1441 2885 -1404
rect 2897 -1444 2921 -1412
rect 2556 -1468 2618 -1444
rect 1716 -1494 1740 -1470
rect 1755 -1480 1789 -1474
rect 1755 -1510 1817 -1480
rect 1783 -1516 1817 -1510
rect 1716 -1549 1740 -1525
rect 2012 -1530 2074 -1506
rect 2186 -1507 2248 -1483
rect 2360 -1503 2422 -1479
rect 1738 -1727 1774 -1687
rect 1780 -1734 1804 -1694
rect 1738 -1836 1774 -1796
rect 1780 -1843 1804 -1803
rect 2084 -1822 2136 -1798
rect 1893 -1851 1930 -1825
rect 1893 -1896 1930 -1870
rect 1739 -1955 1775 -1915
rect 1781 -1962 1805 -1922
rect 1893 -1940 1930 -1914
rect 1893 -1978 1930 -1946
rect 1743 -2063 1779 -2023
rect 1785 -2070 1809 -2030
<< ntransistor >>
rect 2081 -712 2083 -706
rect 2120 -761 2122 -749
rect 2130 -761 2132 -749
rect 2148 -761 2150 -749
rect 2158 -761 2160 -749
rect 2081 -767 2083 -761
rect 2217 -771 2219 -761
rect 2253 -771 2255 -761
rect 2261 -771 2263 -761
rect 2297 -771 2299 -761
rect 2305 -771 2307 -761
rect 2348 -771 2350 -761
rect 2397 -767 2399 -757
rect 2231 -875 2233 -865
rect 2267 -875 2269 -865
rect 2275 -875 2277 -865
rect 2311 -875 2313 -865
rect 2319 -875 2321 -865
rect 2362 -875 2364 -865
rect 2402 -871 2404 -861
rect 931 -893 941 -891
rect 1038 -893 1048 -891
rect 1140 -893 1150 -891
rect 1237 -893 1247 -891
rect 1341 -892 1351 -890
rect 1443 -892 1453 -890
rect 1539 -892 1549 -890
rect 1638 -892 1648 -890
rect 931 -929 941 -927
rect 1038 -929 1048 -927
rect 1140 -929 1150 -927
rect 1237 -929 1247 -927
rect 1341 -928 1351 -926
rect 1443 -928 1453 -926
rect 1539 -928 1549 -926
rect 1638 -928 1648 -926
rect 931 -937 941 -935
rect 1038 -937 1048 -935
rect 1140 -937 1150 -935
rect 1237 -937 1247 -935
rect 1341 -936 1351 -934
rect 1443 -936 1453 -934
rect 1539 -936 1549 -934
rect 1638 -936 1648 -934
rect 2152 -953 2164 -951
rect 2152 -963 2164 -961
rect 931 -973 941 -971
rect 1038 -973 1048 -971
rect 1140 -973 1150 -971
rect 1237 -973 1247 -971
rect 1341 -972 1351 -970
rect 1443 -972 1453 -970
rect 1539 -972 1549 -970
rect 1638 -972 1648 -970
rect 931 -981 941 -979
rect 1038 -981 1048 -979
rect 1140 -981 1150 -979
rect 1237 -981 1247 -979
rect 1341 -980 1351 -978
rect 1443 -980 1453 -978
rect 1539 -980 1549 -978
rect 1638 -980 1648 -978
rect 2152 -981 2164 -979
rect 2152 -991 2164 -989
rect 2321 -1001 2333 -999
rect 2384 -1004 2386 -994
rect 2420 -1004 2422 -994
rect 2428 -1004 2430 -994
rect 2464 -1004 2466 -994
rect 2472 -1004 2474 -994
rect 2515 -1004 2517 -994
rect 2563 -1000 2565 -990
rect 2321 -1011 2333 -1009
rect 931 -1024 941 -1022
rect 1038 -1024 1048 -1022
rect 1140 -1024 1150 -1022
rect 1237 -1024 1247 -1022
rect 1341 -1023 1351 -1021
rect 1443 -1023 1453 -1021
rect 1539 -1023 1549 -1021
rect 1638 -1023 1648 -1021
rect 2109 -1030 2115 -1028
rect 2164 -1030 2170 -1028
rect 2321 -1029 2333 -1027
rect 2321 -1039 2333 -1037
rect 2278 -1078 2284 -1076
rect 2333 -1078 2339 -1076
rect 1716 -1107 1718 -1101
rect 1755 -1156 1757 -1144
rect 1765 -1156 1767 -1144
rect 1783 -1156 1785 -1144
rect 1793 -1156 1795 -1144
rect 1716 -1162 1718 -1156
rect 2504 -1159 2516 -1157
rect 2578 -1162 2580 -1152
rect 2614 -1162 2616 -1152
rect 2622 -1162 2624 -1152
rect 2658 -1162 2660 -1152
rect 2666 -1162 2668 -1152
rect 2709 -1162 2711 -1152
rect 2756 -1158 2758 -1148
rect 2504 -1169 2516 -1167
rect 2504 -1187 2516 -1185
rect 2504 -1197 2516 -1195
rect 1717 -1239 1719 -1233
rect 2461 -1236 2467 -1234
rect 2516 -1236 2522 -1234
rect 2114 -1252 2134 -1250
rect 1756 -1288 1758 -1276
rect 1766 -1288 1768 -1276
rect 1784 -1288 1786 -1276
rect 1794 -1288 1796 -1276
rect 1717 -1294 1719 -1288
rect 2281 -1295 2301 -1293
rect 2463 -1302 2483 -1300
rect 1720 -1383 1722 -1377
rect 1759 -1432 1761 -1420
rect 1769 -1432 1771 -1420
rect 1787 -1432 1789 -1420
rect 1797 -1432 1799 -1420
rect 1720 -1438 1722 -1432
rect 2696 -1469 2698 -1449
rect 2739 -1467 2741 -1457
rect 2775 -1467 2777 -1457
rect 2783 -1467 2785 -1457
rect 2819 -1467 2821 -1457
rect 2827 -1467 2829 -1457
rect 2870 -1467 2872 -1457
rect 2908 -1466 2910 -1456
rect 1727 -1508 1729 -1502
rect 2538 -1542 2638 -1540
rect 1766 -1557 1768 -1545
rect 1776 -1557 1778 -1545
rect 1794 -1557 1796 -1545
rect 1804 -1557 1806 -1545
rect 2350 -1550 2450 -1548
rect 1727 -1563 1729 -1557
rect 2169 -1560 2269 -1558
rect 2001 -1568 2101 -1566
rect 2540 -1651 2640 -1649
rect 2348 -1661 2448 -1659
rect 2168 -1671 2268 -1669
rect 1749 -1770 1751 -1750
rect 1760 -1770 1762 -1750
rect 1791 -1752 1793 -1742
rect 1953 -1779 1955 -1679
rect 2000 -1682 2100 -1680
rect 2033 -1780 2133 -1778
rect 2148 -1811 2168 -1809
rect 1946 -1840 1956 -1838
rect 1749 -1879 1751 -1859
rect 1760 -1879 1762 -1859
rect 1791 -1861 1793 -1851
rect 1946 -1883 1956 -1881
rect 1946 -1891 1956 -1889
rect 1946 -1927 1956 -1925
rect 1946 -1935 1956 -1933
rect 1750 -1998 1752 -1978
rect 1761 -1998 1763 -1978
rect 1792 -1980 1794 -1970
rect 1946 -1971 1956 -1969
rect 1754 -2106 1756 -2086
rect 1765 -2106 1767 -2086
rect 1796 -2088 1798 -2078
<< ptransistor >>
rect 2081 -692 2083 -680
rect 2120 -708 2122 -684
rect 2130 -708 2132 -684
rect 2148 -714 2150 -690
rect 2158 -714 2160 -690
rect 2081 -747 2083 -735
rect 2221 -739 2223 -714
rect 2229 -739 2231 -714
rect 2259 -739 2261 -714
rect 2303 -739 2305 -714
rect 2348 -739 2350 -714
rect 2397 -739 2399 -719
rect 2235 -843 2237 -818
rect 2243 -843 2245 -818
rect 2273 -843 2275 -818
rect 2317 -843 2319 -818
rect 2362 -843 2364 -818
rect 2402 -843 2404 -823
rect 963 -897 988 -895
rect 1070 -897 1095 -895
rect 1172 -897 1197 -895
rect 1269 -897 1294 -895
rect 1373 -896 1398 -894
rect 1475 -896 1500 -894
rect 1571 -896 1596 -894
rect 1670 -896 1695 -894
rect 963 -905 988 -903
rect 1070 -905 1095 -903
rect 1172 -905 1197 -903
rect 1269 -905 1294 -903
rect 1373 -904 1398 -902
rect 1475 -904 1500 -902
rect 1571 -904 1596 -902
rect 1670 -904 1695 -902
rect 963 -935 988 -933
rect 1070 -935 1095 -933
rect 1172 -935 1197 -933
rect 1269 -935 1294 -933
rect 1373 -934 1398 -932
rect 1475 -934 1500 -932
rect 1571 -934 1596 -932
rect 1670 -934 1695 -932
rect 2093 -953 2117 -951
rect 2093 -963 2117 -961
rect 963 -979 988 -977
rect 1070 -979 1095 -977
rect 1172 -979 1197 -977
rect 1269 -979 1294 -977
rect 1373 -978 1398 -976
rect 1475 -978 1500 -976
rect 1571 -978 1596 -976
rect 2388 -972 2390 -947
rect 2396 -972 2398 -947
rect 2426 -972 2428 -947
rect 2470 -972 2472 -947
rect 2515 -972 2517 -947
rect 2563 -972 2565 -952
rect 1670 -978 1695 -976
rect 2087 -981 2111 -979
rect 2087 -991 2111 -989
rect 2262 -1001 2286 -999
rect 2262 -1011 2286 -1009
rect 963 -1024 988 -1022
rect 1070 -1024 1095 -1022
rect 1172 -1024 1197 -1022
rect 1269 -1024 1294 -1022
rect 1373 -1023 1398 -1021
rect 1475 -1023 1500 -1021
rect 1571 -1023 1596 -1021
rect 1670 -1023 1695 -1021
rect 2083 -1030 2095 -1028
rect 2138 -1030 2150 -1028
rect 2256 -1029 2280 -1027
rect 2256 -1039 2280 -1037
rect 1716 -1087 1718 -1075
rect 2252 -1078 2264 -1076
rect 2307 -1078 2319 -1076
rect 1755 -1103 1757 -1079
rect 1765 -1103 1767 -1079
rect 1783 -1109 1785 -1085
rect 1793 -1109 1795 -1085
rect 1716 -1142 1718 -1130
rect 2582 -1130 2584 -1105
rect 2590 -1130 2592 -1105
rect 2620 -1130 2622 -1105
rect 2664 -1130 2666 -1105
rect 2709 -1130 2711 -1105
rect 2756 -1130 2758 -1110
rect 2445 -1159 2469 -1157
rect 2445 -1169 2469 -1167
rect 2439 -1187 2463 -1185
rect 2439 -1197 2463 -1195
rect 1717 -1219 1719 -1207
rect 1756 -1235 1758 -1211
rect 1766 -1235 1768 -1211
rect 1784 -1241 1786 -1217
rect 1794 -1241 1796 -1217
rect 2435 -1236 2447 -1234
rect 2490 -1236 2502 -1234
rect 1717 -1274 1719 -1262
rect 2056 -1252 2096 -1250
rect 2223 -1295 2263 -1293
rect 2405 -1302 2445 -1300
rect 1720 -1363 1722 -1351
rect 1759 -1379 1761 -1355
rect 1769 -1379 1771 -1355
rect 1787 -1385 1789 -1361
rect 1797 -1385 1799 -1361
rect 1720 -1418 1722 -1406
rect 2696 -1431 2698 -1391
rect 2743 -1435 2745 -1410
rect 2751 -1435 2753 -1410
rect 2781 -1435 2783 -1410
rect 2825 -1435 2827 -1410
rect 2870 -1435 2872 -1410
rect 2562 -1457 2612 -1455
rect 2908 -1438 2910 -1418
rect 1727 -1488 1729 -1476
rect 1766 -1504 1768 -1480
rect 1776 -1504 1778 -1480
rect 1794 -1510 1796 -1486
rect 1804 -1510 1806 -1486
rect 2366 -1492 2416 -1490
rect 2192 -1496 2242 -1494
rect 1727 -1543 1729 -1531
rect 2018 -1519 2068 -1517
rect 1749 -1721 1751 -1701
rect 1760 -1721 1762 -1701
rect 1791 -1728 1793 -1708
rect 1749 -1830 1751 -1810
rect 1760 -1830 1762 -1810
rect 2090 -1811 2130 -1809
rect 1791 -1837 1793 -1817
rect 1899 -1840 1924 -1838
rect 1899 -1885 1924 -1883
rect 1899 -1929 1924 -1927
rect 1750 -1949 1752 -1929
rect 1761 -1949 1763 -1929
rect 1792 -1956 1794 -1936
rect 1899 -1959 1924 -1957
rect 1899 -1967 1924 -1965
rect 1754 -2057 1756 -2037
rect 1765 -2057 1767 -2037
rect 1796 -2064 1798 -2044
<< ndiffusion >>
rect 2080 -712 2081 -706
rect 2083 -712 2084 -706
rect 2119 -761 2120 -749
rect 2122 -761 2130 -749
rect 2132 -761 2133 -749
rect 2147 -761 2148 -749
rect 2150 -761 2158 -749
rect 2160 -761 2161 -749
rect 2080 -767 2081 -761
rect 2083 -767 2084 -761
rect 2216 -771 2217 -761
rect 2219 -771 2220 -761
rect 2252 -771 2253 -761
rect 2255 -771 2256 -761
rect 2260 -771 2261 -761
rect 2263 -771 2264 -761
rect 2296 -771 2297 -761
rect 2299 -771 2300 -761
rect 2304 -771 2305 -761
rect 2307 -771 2308 -761
rect 2347 -771 2348 -761
rect 2350 -771 2351 -761
rect 2396 -767 2397 -757
rect 2399 -767 2400 -757
rect 2230 -875 2231 -865
rect 2233 -875 2234 -865
rect 2266 -875 2267 -865
rect 2269 -875 2270 -865
rect 2274 -875 2275 -865
rect 2277 -875 2278 -865
rect 2310 -875 2311 -865
rect 2313 -875 2314 -865
rect 2318 -875 2319 -865
rect 2321 -875 2322 -865
rect 2361 -875 2362 -865
rect 2364 -875 2365 -865
rect 2401 -871 2402 -861
rect 2404 -871 2405 -861
rect 931 -891 941 -890
rect 931 -894 941 -893
rect 1038 -891 1048 -890
rect 1038 -894 1048 -893
rect 1140 -891 1150 -890
rect 1140 -894 1150 -893
rect 1237 -891 1247 -890
rect 1341 -890 1351 -889
rect 1237 -894 1247 -893
rect 1341 -893 1351 -892
rect 1443 -890 1453 -889
rect 1443 -893 1453 -892
rect 1539 -890 1549 -889
rect 1539 -893 1549 -892
rect 1638 -890 1648 -889
rect 1638 -893 1648 -892
rect 931 -927 941 -926
rect 1038 -927 1048 -926
rect 1140 -927 1150 -926
rect 1237 -927 1247 -926
rect 1341 -926 1351 -925
rect 1443 -926 1453 -925
rect 1539 -926 1549 -925
rect 1638 -926 1648 -925
rect 931 -930 941 -929
rect 931 -935 941 -934
rect 1038 -930 1048 -929
rect 1038 -935 1048 -934
rect 1140 -930 1150 -929
rect 1140 -935 1150 -934
rect 1237 -930 1247 -929
rect 1237 -935 1247 -934
rect 1341 -929 1351 -928
rect 1341 -934 1351 -933
rect 1443 -929 1453 -928
rect 1443 -934 1453 -933
rect 1539 -929 1549 -928
rect 1539 -934 1549 -933
rect 1638 -929 1648 -928
rect 1638 -934 1648 -933
rect 931 -938 941 -937
rect 1038 -938 1048 -937
rect 1140 -938 1150 -937
rect 1237 -938 1247 -937
rect 1341 -937 1351 -936
rect 1443 -937 1453 -936
rect 1539 -937 1549 -936
rect 1638 -937 1648 -936
rect 2152 -951 2164 -950
rect 2152 -961 2164 -953
rect 931 -971 941 -970
rect 1038 -971 1048 -970
rect 1140 -971 1150 -970
rect 1237 -971 1247 -970
rect 1341 -970 1351 -969
rect 1443 -970 1453 -969
rect 1539 -970 1549 -969
rect 1638 -970 1648 -969
rect 2152 -964 2164 -963
rect 931 -974 941 -973
rect 931 -979 941 -978
rect 1038 -974 1048 -973
rect 1038 -979 1048 -978
rect 1140 -974 1150 -973
rect 1140 -979 1150 -978
rect 1237 -974 1247 -973
rect 1237 -979 1247 -978
rect 1341 -973 1351 -972
rect 1341 -978 1351 -977
rect 1443 -973 1453 -972
rect 1443 -978 1453 -977
rect 1539 -973 1549 -972
rect 1539 -978 1549 -977
rect 1638 -973 1648 -972
rect 1638 -978 1648 -977
rect 931 -982 941 -981
rect 1038 -982 1048 -981
rect 1140 -982 1150 -981
rect 1237 -982 1247 -981
rect 1341 -981 1351 -980
rect 1443 -981 1453 -980
rect 1539 -981 1549 -980
rect 2152 -979 2164 -978
rect 1638 -981 1648 -980
rect 2152 -989 2164 -981
rect 2152 -992 2164 -991
rect 2321 -999 2333 -998
rect 2321 -1009 2333 -1001
rect 2383 -1004 2384 -994
rect 2386 -1004 2387 -994
rect 2419 -1004 2420 -994
rect 2422 -1004 2423 -994
rect 2427 -1004 2428 -994
rect 2430 -1004 2431 -994
rect 2463 -1004 2464 -994
rect 2466 -1004 2467 -994
rect 2471 -1004 2472 -994
rect 2474 -1004 2475 -994
rect 2514 -1004 2515 -994
rect 2517 -1004 2518 -994
rect 2562 -1000 2563 -990
rect 2565 -1000 2566 -990
rect 2321 -1012 2333 -1011
rect 931 -1022 941 -1021
rect 1038 -1022 1048 -1021
rect 1140 -1022 1150 -1021
rect 1237 -1022 1247 -1021
rect 1341 -1021 1351 -1020
rect 1443 -1021 1453 -1020
rect 1539 -1021 1549 -1020
rect 1638 -1021 1648 -1020
rect 1341 -1024 1351 -1023
rect 931 -1025 941 -1024
rect 1038 -1025 1048 -1024
rect 1140 -1025 1150 -1024
rect 1237 -1025 1247 -1024
rect 1443 -1024 1453 -1023
rect 1539 -1024 1549 -1023
rect 1638 -1024 1648 -1023
rect 2109 -1028 2115 -1027
rect 2321 -1027 2333 -1026
rect 2164 -1028 2170 -1027
rect 2109 -1031 2115 -1030
rect 2164 -1031 2170 -1030
rect 2321 -1037 2333 -1029
rect 2321 -1040 2333 -1039
rect 2278 -1076 2284 -1075
rect 2333 -1076 2339 -1075
rect 1715 -1107 1716 -1101
rect 1718 -1107 1719 -1101
rect 2278 -1079 2284 -1078
rect 2333 -1079 2339 -1078
rect 1754 -1156 1755 -1144
rect 1757 -1156 1765 -1144
rect 1767 -1156 1768 -1144
rect 1782 -1156 1783 -1144
rect 1785 -1156 1793 -1144
rect 1795 -1156 1796 -1144
rect 1715 -1162 1716 -1156
rect 1718 -1162 1719 -1156
rect 2504 -1157 2516 -1156
rect 2504 -1167 2516 -1159
rect 2577 -1162 2578 -1152
rect 2580 -1162 2581 -1152
rect 2613 -1162 2614 -1152
rect 2616 -1162 2617 -1152
rect 2621 -1162 2622 -1152
rect 2624 -1162 2625 -1152
rect 2657 -1162 2658 -1152
rect 2660 -1162 2661 -1152
rect 2665 -1162 2666 -1152
rect 2668 -1162 2669 -1152
rect 2708 -1162 2709 -1152
rect 2711 -1162 2712 -1152
rect 2755 -1158 2756 -1148
rect 2758 -1158 2759 -1148
rect 2504 -1170 2516 -1169
rect 2504 -1185 2516 -1184
rect 2504 -1195 2516 -1187
rect 2504 -1198 2516 -1197
rect 1716 -1239 1717 -1233
rect 1719 -1239 1720 -1233
rect 2461 -1234 2467 -1233
rect 2516 -1234 2522 -1233
rect 2461 -1237 2467 -1236
rect 2516 -1237 2522 -1236
rect 2114 -1250 2134 -1249
rect 2114 -1253 2134 -1252
rect 1755 -1288 1756 -1276
rect 1758 -1288 1766 -1276
rect 1768 -1288 1769 -1276
rect 1783 -1288 1784 -1276
rect 1786 -1288 1794 -1276
rect 1796 -1288 1797 -1276
rect 1716 -1294 1717 -1288
rect 1719 -1294 1720 -1288
rect 2281 -1293 2301 -1292
rect 2281 -1296 2301 -1295
rect 2463 -1300 2483 -1299
rect 2463 -1303 2483 -1302
rect 1719 -1383 1720 -1377
rect 1722 -1383 1723 -1377
rect 1758 -1432 1759 -1420
rect 1761 -1432 1769 -1420
rect 1771 -1432 1772 -1420
rect 1786 -1432 1787 -1420
rect 1789 -1432 1797 -1420
rect 1799 -1432 1800 -1420
rect 1719 -1438 1720 -1432
rect 1722 -1438 1723 -1432
rect 2695 -1469 2696 -1449
rect 2698 -1469 2699 -1449
rect 2738 -1467 2739 -1457
rect 2741 -1467 2742 -1457
rect 2774 -1467 2775 -1457
rect 2777 -1467 2778 -1457
rect 2782 -1467 2783 -1457
rect 2785 -1467 2786 -1457
rect 2818 -1467 2819 -1457
rect 2821 -1467 2822 -1457
rect 2826 -1467 2827 -1457
rect 2829 -1467 2830 -1457
rect 2869 -1467 2870 -1457
rect 2872 -1467 2873 -1457
rect 2907 -1466 2908 -1456
rect 2910 -1466 2911 -1456
rect 1726 -1508 1727 -1502
rect 1729 -1508 1730 -1502
rect 2538 -1540 2638 -1539
rect 2538 -1543 2638 -1542
rect 1765 -1557 1766 -1545
rect 1768 -1557 1776 -1545
rect 1778 -1557 1779 -1545
rect 1793 -1557 1794 -1545
rect 1796 -1557 1804 -1545
rect 1806 -1557 1807 -1545
rect 2350 -1548 2450 -1547
rect 2350 -1551 2450 -1550
rect 1726 -1563 1727 -1557
rect 1729 -1563 1730 -1557
rect 2169 -1558 2269 -1557
rect 2169 -1561 2269 -1560
rect 2001 -1566 2101 -1565
rect 2001 -1569 2101 -1568
rect 2540 -1649 2640 -1648
rect 2540 -1652 2640 -1651
rect 2348 -1659 2448 -1658
rect 2348 -1662 2448 -1661
rect 2168 -1669 2268 -1668
rect 2168 -1672 2268 -1671
rect 1748 -1770 1749 -1750
rect 1751 -1770 1760 -1750
rect 1762 -1770 1763 -1750
rect 1790 -1752 1791 -1742
rect 1793 -1752 1794 -1742
rect 1952 -1779 1953 -1679
rect 1955 -1779 1956 -1679
rect 2000 -1680 2100 -1679
rect 2000 -1683 2100 -1682
rect 2033 -1778 2133 -1777
rect 2033 -1781 2133 -1780
rect 2148 -1809 2168 -1808
rect 2148 -1812 2168 -1811
rect 1946 -1838 1956 -1837
rect 1946 -1841 1956 -1840
rect 1748 -1879 1749 -1859
rect 1751 -1879 1760 -1859
rect 1762 -1879 1763 -1859
rect 1790 -1861 1791 -1851
rect 1793 -1861 1794 -1851
rect 1946 -1881 1956 -1880
rect 1946 -1884 1956 -1883
rect 1946 -1889 1956 -1888
rect 1946 -1892 1956 -1891
rect 1946 -1925 1956 -1924
rect 1946 -1928 1956 -1927
rect 1946 -1933 1956 -1932
rect 1946 -1936 1956 -1935
rect 1749 -1998 1750 -1978
rect 1752 -1998 1761 -1978
rect 1763 -1998 1764 -1978
rect 1791 -1980 1792 -1970
rect 1794 -1980 1795 -1970
rect 1946 -1969 1956 -1968
rect 1946 -1972 1956 -1971
rect 1753 -2106 1754 -2086
rect 1756 -2106 1765 -2086
rect 1767 -2106 1768 -2086
rect 1795 -2088 1796 -2078
rect 1798 -2088 1799 -2078
<< pdiffusion >>
rect 2080 -692 2081 -680
rect 2083 -692 2084 -680
rect 2119 -708 2120 -684
rect 2122 -708 2124 -684
rect 2128 -708 2130 -684
rect 2132 -708 2133 -684
rect 2147 -714 2148 -690
rect 2150 -714 2152 -690
rect 2156 -714 2158 -690
rect 2160 -714 2161 -690
rect 2080 -747 2081 -735
rect 2083 -747 2084 -735
rect 2220 -739 2221 -714
rect 2223 -739 2224 -714
rect 2228 -739 2229 -714
rect 2231 -739 2232 -714
rect 2258 -739 2259 -714
rect 2261 -739 2262 -714
rect 2302 -739 2303 -714
rect 2305 -739 2306 -714
rect 2347 -739 2348 -714
rect 2350 -739 2351 -714
rect 2396 -739 2397 -719
rect 2399 -739 2400 -719
rect 2234 -843 2235 -818
rect 2237 -843 2238 -818
rect 2242 -843 2243 -818
rect 2245 -843 2246 -818
rect 2272 -843 2273 -818
rect 2275 -843 2276 -818
rect 2316 -843 2317 -818
rect 2319 -843 2320 -818
rect 2361 -843 2362 -818
rect 2364 -843 2365 -818
rect 2401 -843 2402 -823
rect 2404 -843 2405 -823
rect 963 -895 988 -894
rect 963 -898 988 -897
rect 1070 -895 1095 -894
rect 1070 -898 1095 -897
rect 1172 -895 1197 -894
rect 1172 -898 1197 -897
rect 1269 -895 1294 -894
rect 1373 -894 1398 -893
rect 1373 -897 1398 -896
rect 1475 -894 1500 -893
rect 1475 -897 1500 -896
rect 1571 -894 1596 -893
rect 1571 -897 1596 -896
rect 1670 -894 1695 -893
rect 1670 -897 1695 -896
rect 1269 -898 1294 -897
rect 963 -903 988 -902
rect 1070 -903 1095 -902
rect 1172 -903 1197 -902
rect 1269 -903 1294 -902
rect 1373 -902 1398 -901
rect 1475 -902 1500 -901
rect 1571 -902 1596 -901
rect 1670 -902 1695 -901
rect 1373 -905 1398 -904
rect 963 -906 988 -905
rect 1070 -906 1095 -905
rect 1172 -906 1197 -905
rect 1269 -906 1294 -905
rect 1475 -905 1500 -904
rect 1571 -905 1596 -904
rect 1670 -905 1695 -904
rect 963 -933 988 -932
rect 1070 -933 1095 -932
rect 1172 -933 1197 -932
rect 1269 -933 1294 -932
rect 1373 -932 1398 -931
rect 1475 -932 1500 -931
rect 1571 -932 1596 -931
rect 1670 -932 1695 -931
rect 963 -936 988 -935
rect 1070 -936 1095 -935
rect 1172 -936 1197 -935
rect 1269 -936 1294 -935
rect 1373 -935 1398 -934
rect 1475 -935 1500 -934
rect 1571 -935 1596 -934
rect 1670 -935 1695 -934
rect 2093 -951 2117 -950
rect 2093 -955 2117 -953
rect 2093 -961 2117 -959
rect 2093 -964 2117 -963
rect 963 -977 988 -976
rect 1070 -977 1095 -976
rect 1172 -977 1197 -976
rect 1269 -977 1294 -976
rect 1373 -976 1398 -975
rect 1475 -976 1500 -975
rect 1571 -976 1596 -975
rect 2387 -972 2388 -947
rect 2390 -972 2391 -947
rect 2395 -972 2396 -947
rect 2398 -972 2399 -947
rect 2425 -972 2426 -947
rect 2428 -972 2429 -947
rect 2469 -972 2470 -947
rect 2472 -972 2473 -947
rect 2514 -972 2515 -947
rect 2517 -972 2518 -947
rect 2562 -972 2563 -952
rect 2565 -972 2566 -952
rect 1670 -976 1695 -975
rect 963 -980 988 -979
rect 1070 -980 1095 -979
rect 1172 -980 1197 -979
rect 1269 -980 1294 -979
rect 1373 -979 1398 -978
rect 1475 -979 1500 -978
rect 1571 -979 1596 -978
rect 1670 -979 1695 -978
rect 2087 -979 2111 -978
rect 2087 -983 2111 -981
rect 2087 -989 2111 -987
rect 2087 -992 2111 -991
rect 2262 -999 2286 -998
rect 2262 -1003 2286 -1001
rect 2262 -1009 2286 -1007
rect 2262 -1012 2286 -1011
rect 963 -1022 988 -1021
rect 1070 -1022 1095 -1021
rect 1172 -1022 1197 -1021
rect 1373 -1021 1398 -1020
rect 1475 -1021 1500 -1020
rect 1571 -1021 1596 -1020
rect 1670 -1021 1695 -1020
rect 1269 -1022 1294 -1021
rect 963 -1025 988 -1024
rect 1070 -1025 1095 -1024
rect 1172 -1025 1197 -1024
rect 1269 -1025 1294 -1024
rect 1373 -1024 1398 -1023
rect 1475 -1024 1500 -1023
rect 1571 -1024 1596 -1023
rect 1670 -1024 1695 -1023
rect 2083 -1028 2095 -1027
rect 2138 -1028 2150 -1027
rect 2256 -1027 2280 -1026
rect 2083 -1031 2095 -1030
rect 2138 -1031 2150 -1030
rect 2256 -1031 2280 -1029
rect 2256 -1037 2280 -1035
rect 2256 -1040 2280 -1039
rect 1715 -1087 1716 -1075
rect 1718 -1087 1719 -1075
rect 2252 -1076 2264 -1075
rect 2307 -1076 2319 -1075
rect 2252 -1079 2264 -1078
rect 1754 -1103 1755 -1079
rect 1757 -1103 1759 -1079
rect 1763 -1103 1765 -1079
rect 1767 -1103 1768 -1079
rect 2307 -1079 2319 -1078
rect 1782 -1109 1783 -1085
rect 1785 -1109 1787 -1085
rect 1791 -1109 1793 -1085
rect 1795 -1109 1796 -1085
rect 1715 -1142 1716 -1130
rect 1718 -1142 1719 -1130
rect 2581 -1130 2582 -1105
rect 2584 -1130 2585 -1105
rect 2589 -1130 2590 -1105
rect 2592 -1130 2593 -1105
rect 2619 -1130 2620 -1105
rect 2622 -1130 2623 -1105
rect 2663 -1130 2664 -1105
rect 2666 -1130 2667 -1105
rect 2708 -1130 2709 -1105
rect 2711 -1130 2712 -1105
rect 2755 -1130 2756 -1110
rect 2758 -1130 2759 -1110
rect 2445 -1157 2469 -1156
rect 2445 -1161 2469 -1159
rect 2445 -1167 2469 -1165
rect 2445 -1170 2469 -1169
rect 2439 -1185 2463 -1184
rect 2439 -1189 2463 -1187
rect 2439 -1195 2463 -1193
rect 2439 -1198 2463 -1197
rect 1716 -1219 1717 -1207
rect 1719 -1219 1720 -1207
rect 1755 -1235 1756 -1211
rect 1758 -1235 1760 -1211
rect 1764 -1235 1766 -1211
rect 1768 -1235 1769 -1211
rect 1783 -1241 1784 -1217
rect 1786 -1241 1788 -1217
rect 1792 -1241 1794 -1217
rect 1796 -1241 1797 -1217
rect 2435 -1234 2447 -1233
rect 2490 -1234 2502 -1233
rect 2435 -1237 2447 -1236
rect 2490 -1237 2502 -1236
rect 1716 -1274 1717 -1262
rect 1719 -1274 1720 -1262
rect 2056 -1250 2096 -1249
rect 2056 -1253 2096 -1252
rect 2223 -1293 2263 -1292
rect 2223 -1296 2263 -1295
rect 2405 -1300 2445 -1299
rect 2405 -1303 2445 -1302
rect 1719 -1363 1720 -1351
rect 1722 -1363 1723 -1351
rect 1758 -1379 1759 -1355
rect 1761 -1379 1763 -1355
rect 1767 -1379 1769 -1355
rect 1771 -1379 1772 -1355
rect 1786 -1385 1787 -1361
rect 1789 -1385 1791 -1361
rect 1795 -1385 1797 -1361
rect 1799 -1385 1800 -1361
rect 1719 -1418 1720 -1406
rect 1722 -1418 1723 -1406
rect 2695 -1431 2696 -1391
rect 2698 -1431 2699 -1391
rect 2742 -1435 2743 -1410
rect 2745 -1435 2746 -1410
rect 2750 -1435 2751 -1410
rect 2753 -1435 2754 -1410
rect 2780 -1435 2781 -1410
rect 2783 -1435 2784 -1410
rect 2824 -1435 2825 -1410
rect 2827 -1435 2828 -1410
rect 2869 -1435 2870 -1410
rect 2872 -1435 2873 -1410
rect 2562 -1455 2612 -1454
rect 2562 -1458 2612 -1457
rect 2907 -1438 2908 -1418
rect 2910 -1438 2911 -1418
rect 1726 -1488 1727 -1476
rect 1729 -1488 1730 -1476
rect 1765 -1504 1766 -1480
rect 1768 -1504 1770 -1480
rect 1774 -1504 1776 -1480
rect 1778 -1504 1779 -1480
rect 1793 -1510 1794 -1486
rect 1796 -1510 1798 -1486
rect 1802 -1510 1804 -1486
rect 1806 -1510 1807 -1486
rect 2192 -1494 2242 -1493
rect 2366 -1490 2416 -1489
rect 2366 -1493 2416 -1492
rect 2192 -1497 2242 -1496
rect 1726 -1543 1727 -1531
rect 1729 -1543 1730 -1531
rect 2018 -1517 2068 -1516
rect 2018 -1520 2068 -1519
rect 1748 -1721 1749 -1701
rect 1751 -1721 1755 -1701
rect 1759 -1721 1760 -1701
rect 1762 -1721 1763 -1701
rect 1790 -1728 1791 -1708
rect 1793 -1728 1794 -1708
rect 2090 -1809 2130 -1808
rect 1748 -1830 1749 -1810
rect 1751 -1830 1755 -1810
rect 1759 -1830 1760 -1810
rect 1762 -1830 1763 -1810
rect 2090 -1812 2130 -1811
rect 1790 -1837 1791 -1817
rect 1793 -1837 1794 -1817
rect 1899 -1838 1924 -1837
rect 1899 -1841 1924 -1840
rect 1899 -1883 1924 -1882
rect 1899 -1886 1924 -1885
rect 1899 -1927 1924 -1926
rect 1749 -1949 1750 -1929
rect 1752 -1949 1756 -1929
rect 1760 -1949 1761 -1929
rect 1763 -1949 1764 -1929
rect 1899 -1930 1924 -1929
rect 1791 -1956 1792 -1936
rect 1794 -1956 1795 -1936
rect 1899 -1957 1924 -1956
rect 1899 -1960 1924 -1959
rect 1899 -1965 1924 -1964
rect 1899 -1968 1924 -1967
rect 1753 -2057 1754 -2037
rect 1756 -2057 1760 -2037
rect 1764 -2057 1765 -2037
rect 1767 -2057 1768 -2037
rect 1795 -2064 1796 -2044
rect 1798 -2064 1799 -2044
<< ndcontact >>
rect 2076 -712 2080 -706
rect 2084 -712 2088 -706
rect 2115 -761 2119 -749
rect 2133 -761 2137 -749
rect 2143 -761 2147 -749
rect 2161 -761 2165 -749
rect 2076 -767 2080 -761
rect 2084 -767 2088 -761
rect 2212 -771 2216 -761
rect 2220 -771 2224 -761
rect 2248 -771 2252 -761
rect 2256 -771 2260 -761
rect 2264 -771 2268 -761
rect 2292 -771 2296 -761
rect 2300 -771 2304 -761
rect 2308 -771 2312 -761
rect 2343 -771 2347 -761
rect 2351 -771 2355 -761
rect 2392 -767 2396 -757
rect 2400 -767 2404 -757
rect 2226 -875 2230 -865
rect 2234 -875 2238 -865
rect 2262 -875 2266 -865
rect 2270 -875 2274 -865
rect 2278 -875 2282 -865
rect 2306 -875 2310 -865
rect 2314 -875 2318 -865
rect 2322 -875 2326 -865
rect 2357 -875 2361 -865
rect 2365 -875 2369 -865
rect 2397 -871 2401 -861
rect 2405 -871 2409 -861
rect 931 -890 941 -886
rect 1038 -890 1048 -886
rect 931 -898 941 -894
rect 1140 -890 1150 -886
rect 1038 -898 1048 -894
rect 1237 -890 1247 -886
rect 1140 -898 1150 -894
rect 1341 -889 1351 -885
rect 1443 -889 1453 -885
rect 1237 -898 1247 -894
rect 1341 -897 1351 -893
rect 1539 -889 1549 -885
rect 1443 -897 1453 -893
rect 1638 -889 1648 -885
rect 1539 -897 1549 -893
rect 1638 -897 1648 -893
rect 931 -926 941 -922
rect 1038 -926 1048 -922
rect 1140 -926 1150 -922
rect 1237 -926 1247 -922
rect 1341 -925 1351 -921
rect 1443 -925 1453 -921
rect 1539 -925 1549 -921
rect 1638 -925 1648 -921
rect 931 -934 941 -930
rect 1038 -934 1048 -930
rect 1140 -934 1150 -930
rect 1237 -934 1247 -930
rect 1341 -933 1351 -929
rect 1443 -933 1453 -929
rect 1539 -933 1549 -929
rect 1638 -933 1648 -929
rect 931 -942 941 -938
rect 1038 -942 1048 -938
rect 1140 -942 1150 -938
rect 1237 -942 1247 -938
rect 1341 -941 1351 -937
rect 1443 -941 1453 -937
rect 1539 -941 1549 -937
rect 1638 -941 1648 -937
rect 2152 -950 2164 -946
rect 931 -970 941 -966
rect 1038 -970 1048 -966
rect 1140 -970 1150 -966
rect 1237 -970 1247 -966
rect 1341 -969 1351 -965
rect 1443 -969 1453 -965
rect 1539 -969 1549 -965
rect 1638 -969 1648 -965
rect 2152 -968 2164 -964
rect 931 -978 941 -974
rect 1038 -978 1048 -974
rect 1140 -978 1150 -974
rect 1237 -978 1247 -974
rect 1341 -977 1351 -973
rect 1443 -977 1453 -973
rect 1539 -977 1549 -973
rect 1638 -977 1648 -973
rect 931 -986 941 -982
rect 1038 -986 1048 -982
rect 1140 -986 1150 -982
rect 1237 -986 1247 -982
rect 1341 -985 1351 -981
rect 1443 -985 1453 -981
rect 1539 -985 1549 -981
rect 2152 -978 2164 -974
rect 1638 -985 1648 -981
rect 2152 -996 2164 -992
rect 2321 -998 2333 -994
rect 2379 -1004 2383 -994
rect 2387 -1004 2391 -994
rect 2415 -1004 2419 -994
rect 2423 -1004 2427 -994
rect 2431 -1004 2435 -994
rect 2459 -1004 2463 -994
rect 2467 -1004 2471 -994
rect 2475 -1004 2479 -994
rect 2510 -1004 2514 -994
rect 2518 -1004 2522 -994
rect 2558 -1000 2562 -990
rect 2566 -1000 2570 -990
rect 2321 -1016 2333 -1012
rect 931 -1021 941 -1017
rect 1038 -1021 1048 -1017
rect 1140 -1021 1150 -1017
rect 1237 -1021 1247 -1017
rect 1341 -1020 1351 -1016
rect 1443 -1020 1453 -1016
rect 1539 -1020 1549 -1016
rect 1638 -1020 1648 -1016
rect 931 -1029 941 -1025
rect 1038 -1029 1048 -1025
rect 1140 -1029 1150 -1025
rect 1237 -1029 1247 -1025
rect 1341 -1028 1351 -1024
rect 1443 -1028 1453 -1024
rect 1539 -1028 1549 -1024
rect 1638 -1028 1648 -1024
rect 2109 -1027 2115 -1023
rect 2164 -1027 2170 -1023
rect 2321 -1026 2333 -1022
rect 2109 -1035 2115 -1031
rect 2164 -1035 2170 -1031
rect 2321 -1044 2333 -1040
rect 2278 -1075 2284 -1071
rect 2333 -1075 2339 -1071
rect 1711 -1107 1715 -1101
rect 1719 -1107 1723 -1101
rect 2278 -1083 2284 -1079
rect 2333 -1083 2339 -1079
rect 1750 -1156 1754 -1144
rect 1768 -1156 1772 -1144
rect 1778 -1156 1782 -1144
rect 1796 -1156 1800 -1144
rect 2504 -1156 2516 -1152
rect 1711 -1162 1715 -1156
rect 1719 -1162 1723 -1156
rect 2573 -1162 2577 -1152
rect 2581 -1162 2585 -1152
rect 2609 -1162 2613 -1152
rect 2617 -1162 2621 -1152
rect 2625 -1162 2629 -1152
rect 2653 -1162 2657 -1152
rect 2661 -1162 2665 -1152
rect 2669 -1162 2673 -1152
rect 2704 -1162 2708 -1152
rect 2712 -1162 2716 -1152
rect 2751 -1158 2755 -1148
rect 2759 -1158 2763 -1148
rect 2504 -1174 2516 -1170
rect 2504 -1184 2516 -1180
rect 2504 -1202 2516 -1198
rect 1712 -1239 1716 -1233
rect 1720 -1239 1724 -1233
rect 2461 -1233 2467 -1229
rect 2516 -1233 2522 -1229
rect 2461 -1241 2467 -1237
rect 2516 -1241 2522 -1237
rect 2114 -1249 2134 -1245
rect 2114 -1257 2134 -1253
rect 1751 -1288 1755 -1276
rect 1769 -1288 1773 -1276
rect 1779 -1288 1783 -1276
rect 1797 -1288 1801 -1276
rect 1712 -1294 1716 -1288
rect 1720 -1294 1724 -1288
rect 2281 -1292 2301 -1288
rect 2281 -1300 2301 -1296
rect 2463 -1299 2483 -1295
rect 2463 -1307 2483 -1303
rect 1715 -1383 1719 -1377
rect 1723 -1383 1727 -1377
rect 1754 -1432 1758 -1420
rect 1772 -1432 1776 -1420
rect 1782 -1432 1786 -1420
rect 1800 -1432 1804 -1420
rect 1715 -1438 1719 -1432
rect 1723 -1438 1727 -1432
rect 2691 -1469 2695 -1449
rect 2699 -1469 2703 -1449
rect 2734 -1467 2738 -1457
rect 2742 -1467 2746 -1457
rect 2770 -1467 2774 -1457
rect 2778 -1467 2782 -1457
rect 2786 -1467 2790 -1457
rect 2814 -1467 2818 -1457
rect 2822 -1467 2826 -1457
rect 2830 -1467 2834 -1457
rect 2865 -1467 2869 -1457
rect 2873 -1467 2877 -1457
rect 2903 -1466 2907 -1456
rect 2911 -1466 2915 -1456
rect 1722 -1508 1726 -1502
rect 1730 -1508 1734 -1502
rect 2538 -1539 2638 -1535
rect 1761 -1557 1765 -1545
rect 1779 -1557 1783 -1545
rect 1789 -1557 1793 -1545
rect 1807 -1557 1811 -1545
rect 2350 -1547 2450 -1543
rect 2538 -1547 2638 -1543
rect 1722 -1563 1726 -1557
rect 1730 -1563 1734 -1557
rect 2169 -1557 2269 -1553
rect 2350 -1555 2450 -1551
rect 2001 -1565 2101 -1561
rect 2169 -1565 2269 -1561
rect 2001 -1573 2101 -1569
rect 2540 -1648 2640 -1644
rect 2348 -1658 2448 -1654
rect 2540 -1656 2640 -1652
rect 2168 -1668 2268 -1664
rect 2348 -1666 2448 -1662
rect 1744 -1770 1748 -1750
rect 1763 -1770 1767 -1750
rect 1786 -1752 1790 -1742
rect 1794 -1752 1798 -1742
rect 1948 -1779 1952 -1679
rect 1956 -1779 1960 -1679
rect 2000 -1679 2100 -1675
rect 2168 -1676 2268 -1672
rect 2000 -1687 2100 -1683
rect 2033 -1777 2133 -1773
rect 2033 -1785 2133 -1781
rect 2148 -1808 2168 -1804
rect 2148 -1816 2168 -1812
rect 1946 -1837 1956 -1833
rect 1946 -1845 1956 -1841
rect 1744 -1879 1748 -1859
rect 1763 -1879 1767 -1859
rect 1786 -1861 1790 -1851
rect 1794 -1861 1798 -1851
rect 1946 -1880 1956 -1876
rect 1946 -1888 1956 -1884
rect 1946 -1896 1956 -1892
rect 1946 -1924 1956 -1920
rect 1946 -1932 1956 -1928
rect 1946 -1940 1956 -1936
rect 1745 -1998 1749 -1978
rect 1764 -1998 1768 -1978
rect 1787 -1980 1791 -1970
rect 1795 -1980 1799 -1970
rect 1946 -1968 1956 -1964
rect 1946 -1976 1956 -1972
rect 1749 -2106 1753 -2086
rect 1768 -2106 1772 -2086
rect 1791 -2088 1795 -2078
rect 1799 -2088 1803 -2078
<< pdcontact >>
rect 2076 -692 2080 -680
rect 2084 -692 2088 -680
rect 2115 -708 2119 -684
rect 2124 -708 2128 -684
rect 2133 -708 2137 -684
rect 2143 -714 2147 -690
rect 2152 -714 2156 -690
rect 2161 -714 2165 -690
rect 2076 -747 2080 -735
rect 2084 -747 2088 -735
rect 2216 -739 2220 -714
rect 2224 -739 2228 -714
rect 2232 -739 2236 -714
rect 2254 -739 2258 -714
rect 2262 -739 2266 -714
rect 2298 -739 2302 -714
rect 2306 -739 2310 -714
rect 2343 -739 2347 -714
rect 2351 -739 2355 -714
rect 2392 -739 2396 -719
rect 2400 -739 2404 -719
rect 2230 -843 2234 -818
rect 2238 -843 2242 -818
rect 2246 -843 2250 -818
rect 2268 -843 2272 -818
rect 2276 -843 2280 -818
rect 2312 -843 2316 -818
rect 2320 -843 2324 -818
rect 2357 -843 2361 -818
rect 2365 -843 2369 -818
rect 2397 -843 2401 -823
rect 2405 -843 2409 -823
rect 963 -894 988 -890
rect 1070 -894 1095 -890
rect 1172 -894 1197 -890
rect 1269 -894 1294 -890
rect 1373 -893 1398 -889
rect 1475 -893 1500 -889
rect 1571 -893 1596 -889
rect 1670 -893 1695 -889
rect 963 -902 988 -898
rect 1070 -902 1095 -898
rect 1172 -902 1197 -898
rect 1269 -902 1294 -898
rect 1373 -901 1398 -897
rect 1475 -901 1500 -897
rect 1571 -901 1596 -897
rect 1670 -901 1695 -897
rect 963 -910 988 -906
rect 1070 -910 1095 -906
rect 1172 -910 1197 -906
rect 1269 -910 1294 -906
rect 1373 -909 1398 -905
rect 1475 -909 1500 -905
rect 1571 -909 1596 -905
rect 1670 -909 1695 -905
rect 963 -932 988 -928
rect 1070 -932 1095 -928
rect 1172 -932 1197 -928
rect 1269 -932 1294 -928
rect 1373 -931 1398 -927
rect 1475 -931 1500 -927
rect 1571 -931 1596 -927
rect 1670 -931 1695 -927
rect 963 -940 988 -936
rect 1070 -940 1095 -936
rect 1172 -940 1197 -936
rect 1269 -940 1294 -936
rect 1373 -939 1398 -935
rect 1475 -939 1500 -935
rect 1571 -939 1596 -935
rect 1670 -939 1695 -935
rect 2093 -950 2117 -946
rect 2093 -959 2117 -955
rect 2093 -968 2117 -964
rect 963 -976 988 -972
rect 1070 -976 1095 -972
rect 1172 -976 1197 -972
rect 1269 -976 1294 -972
rect 1373 -975 1398 -971
rect 1475 -975 1500 -971
rect 1571 -975 1596 -971
rect 1670 -975 1695 -971
rect 2383 -972 2387 -947
rect 2391 -972 2395 -947
rect 2399 -972 2403 -947
rect 2421 -972 2425 -947
rect 2429 -972 2433 -947
rect 2465 -972 2469 -947
rect 2473 -972 2477 -947
rect 2510 -972 2514 -947
rect 2518 -972 2522 -947
rect 2558 -972 2562 -952
rect 2566 -972 2570 -952
rect 2087 -978 2111 -974
rect 963 -984 988 -980
rect 1070 -984 1095 -980
rect 1172 -984 1197 -980
rect 1269 -984 1294 -980
rect 1373 -983 1398 -979
rect 1475 -983 1500 -979
rect 1571 -983 1596 -979
rect 1670 -983 1695 -979
rect 2087 -987 2111 -983
rect 2087 -996 2111 -992
rect 2262 -998 2286 -994
rect 2262 -1007 2286 -1003
rect 2262 -1016 2286 -1012
rect 963 -1021 988 -1017
rect 1070 -1021 1095 -1017
rect 1172 -1021 1197 -1017
rect 1269 -1021 1294 -1017
rect 1373 -1020 1398 -1016
rect 1475 -1020 1500 -1016
rect 1571 -1020 1596 -1016
rect 1670 -1020 1695 -1016
rect 963 -1029 988 -1025
rect 1070 -1029 1095 -1025
rect 1172 -1029 1197 -1025
rect 1269 -1029 1294 -1025
rect 1373 -1028 1398 -1024
rect 1475 -1028 1500 -1024
rect 1571 -1028 1596 -1024
rect 1670 -1028 1695 -1024
rect 2083 -1027 2095 -1023
rect 2138 -1027 2150 -1023
rect 2256 -1026 2280 -1022
rect 2083 -1035 2095 -1031
rect 2138 -1035 2150 -1031
rect 2256 -1035 2280 -1031
rect 2256 -1044 2280 -1040
rect 2252 -1075 2264 -1071
rect 1711 -1087 1715 -1075
rect 1719 -1087 1723 -1075
rect 2307 -1075 2319 -1071
rect 1750 -1103 1754 -1079
rect 1759 -1103 1763 -1079
rect 1768 -1103 1772 -1079
rect 2252 -1083 2264 -1079
rect 2307 -1083 2319 -1079
rect 1778 -1109 1782 -1085
rect 1787 -1109 1791 -1085
rect 1796 -1109 1800 -1085
rect 1711 -1142 1715 -1130
rect 1719 -1142 1723 -1130
rect 2577 -1130 2581 -1105
rect 2585 -1130 2589 -1105
rect 2593 -1130 2597 -1105
rect 2615 -1130 2619 -1105
rect 2623 -1130 2627 -1105
rect 2659 -1130 2663 -1105
rect 2667 -1130 2671 -1105
rect 2704 -1130 2708 -1105
rect 2712 -1130 2716 -1105
rect 2751 -1130 2755 -1110
rect 2759 -1130 2763 -1110
rect 2445 -1156 2469 -1152
rect 2445 -1165 2469 -1161
rect 2445 -1174 2469 -1170
rect 2439 -1184 2463 -1180
rect 2439 -1193 2463 -1189
rect 2439 -1202 2463 -1198
rect 1712 -1219 1716 -1207
rect 1720 -1219 1724 -1207
rect 1751 -1235 1755 -1211
rect 1760 -1235 1764 -1211
rect 1769 -1235 1773 -1211
rect 1779 -1241 1783 -1217
rect 1788 -1241 1792 -1217
rect 1797 -1241 1801 -1217
rect 2435 -1233 2447 -1229
rect 2490 -1233 2502 -1229
rect 2435 -1241 2447 -1237
rect 2490 -1241 2502 -1237
rect 1712 -1274 1716 -1262
rect 1720 -1274 1724 -1262
rect 2056 -1249 2096 -1245
rect 2056 -1257 2096 -1253
rect 2223 -1292 2263 -1288
rect 2223 -1300 2263 -1296
rect 2405 -1299 2445 -1295
rect 2405 -1307 2445 -1303
rect 1715 -1363 1719 -1351
rect 1723 -1363 1727 -1351
rect 1754 -1379 1758 -1355
rect 1763 -1379 1767 -1355
rect 1772 -1379 1776 -1355
rect 1782 -1385 1786 -1361
rect 1791 -1385 1795 -1361
rect 1800 -1385 1804 -1361
rect 1715 -1418 1719 -1406
rect 1723 -1418 1727 -1406
rect 2691 -1431 2695 -1391
rect 2699 -1431 2703 -1391
rect 2738 -1435 2742 -1410
rect 2746 -1435 2750 -1410
rect 2754 -1435 2758 -1410
rect 2776 -1435 2780 -1410
rect 2784 -1435 2788 -1410
rect 2820 -1435 2824 -1410
rect 2828 -1435 2832 -1410
rect 2865 -1435 2869 -1410
rect 2873 -1435 2877 -1410
rect 2562 -1454 2612 -1450
rect 2562 -1462 2612 -1458
rect 2903 -1438 2907 -1418
rect 2911 -1438 2915 -1418
rect 1722 -1488 1726 -1476
rect 1730 -1488 1734 -1476
rect 1761 -1504 1765 -1480
rect 1770 -1504 1774 -1480
rect 1779 -1504 1783 -1480
rect 1789 -1510 1793 -1486
rect 1798 -1510 1802 -1486
rect 1807 -1510 1811 -1486
rect 2192 -1493 2242 -1489
rect 2366 -1489 2416 -1485
rect 2366 -1497 2416 -1493
rect 2192 -1501 2242 -1497
rect 1722 -1543 1726 -1531
rect 1730 -1543 1734 -1531
rect 2018 -1516 2068 -1512
rect 2018 -1524 2068 -1520
rect 1744 -1721 1748 -1701
rect 1755 -1721 1759 -1701
rect 1763 -1721 1767 -1701
rect 1786 -1728 1790 -1708
rect 1794 -1728 1798 -1708
rect 2090 -1808 2130 -1804
rect 1744 -1830 1748 -1810
rect 1755 -1830 1759 -1810
rect 1763 -1830 1767 -1810
rect 2090 -1816 2130 -1812
rect 1786 -1837 1790 -1817
rect 1794 -1837 1798 -1817
rect 1899 -1837 1924 -1833
rect 1899 -1845 1924 -1841
rect 1899 -1882 1924 -1878
rect 1899 -1890 1924 -1886
rect 1899 -1926 1924 -1922
rect 1745 -1949 1749 -1929
rect 1756 -1949 1760 -1929
rect 1764 -1949 1768 -1929
rect 1899 -1934 1924 -1930
rect 1787 -1956 1791 -1936
rect 1795 -1956 1799 -1936
rect 1899 -1956 1924 -1952
rect 1899 -1964 1924 -1960
rect 1899 -1972 1924 -1968
rect 1749 -2057 1753 -2037
rect 1760 -2057 1764 -2037
rect 1768 -2057 1772 -2037
rect 1791 -2064 1795 -2044
rect 1799 -2064 1803 -2044
<< psubstratepcontact >>
rect 1800 -1761 1805 -1757
rect 1800 -1870 1805 -1866
rect 1801 -1989 1806 -1985
rect 1805 -2097 1810 -2093
<< nsubstratencontact >>
rect 2387 -713 2391 -709
rect 2392 -817 2396 -813
rect 2553 -946 2557 -942
rect 2746 -1104 2750 -1100
rect 2046 -1262 2050 -1258
rect 2213 -1305 2217 -1301
rect 2395 -1312 2399 -1308
rect 2686 -1385 2690 -1381
rect 2551 -1449 2556 -1445
rect 2898 -1412 2902 -1408
rect 2355 -1484 2360 -1480
rect 2181 -1488 2186 -1484
rect 2007 -1511 2012 -1507
rect 1744 -1696 1748 -1690
rect 1796 -1701 1800 -1697
rect 1744 -1805 1748 -1799
rect 1796 -1810 1800 -1806
rect 2080 -1821 2084 -1817
rect 1745 -1924 1749 -1918
rect 1797 -1929 1801 -1925
rect 1749 -2032 1753 -2026
rect 1801 -2037 1805 -2033
<< polysilicon >>
rect 2081 -680 2083 -677
rect 2120 -684 2122 -681
rect 2130 -684 2132 -681
rect 2081 -706 2083 -692
rect 2148 -690 2150 -687
rect 2158 -690 2160 -687
rect 2081 -715 2083 -712
rect 2120 -717 2122 -708
rect 2130 -718 2132 -708
rect 2221 -714 2223 -711
rect 2229 -714 2231 -711
rect 2259 -714 2261 -711
rect 2303 -714 2305 -711
rect 2348 -714 2350 -711
rect 2081 -735 2083 -732
rect 2081 -761 2083 -747
rect 2120 -749 2122 -722
rect 2130 -749 2132 -723
rect 2148 -725 2150 -714
rect 2148 -749 2150 -729
rect 2158 -736 2160 -714
rect 2397 -719 2399 -716
rect 2158 -749 2160 -740
rect 2221 -746 2223 -739
rect 2216 -750 2223 -746
rect 2217 -761 2219 -750
rect 2229 -758 2231 -739
rect 2259 -747 2261 -739
rect 2303 -747 2305 -739
rect 2253 -749 2261 -747
rect 2297 -749 2305 -747
rect 2253 -761 2255 -749
rect 2261 -761 2263 -752
rect 2297 -761 2299 -749
rect 2305 -761 2307 -752
rect 2348 -761 2350 -739
rect 2397 -757 2399 -739
rect 2120 -764 2122 -761
rect 2130 -764 2132 -761
rect 2148 -764 2150 -761
rect 2158 -764 2160 -761
rect 2081 -770 2083 -767
rect 2397 -771 2399 -767
rect 2217 -774 2219 -771
rect 2253 -774 2255 -771
rect 2261 -774 2263 -771
rect 2297 -774 2299 -771
rect 2305 -774 2307 -771
rect 2348 -774 2350 -771
rect 2235 -818 2237 -815
rect 2243 -818 2245 -815
rect 2273 -818 2275 -815
rect 2317 -818 2319 -815
rect 2362 -818 2364 -815
rect 2402 -823 2404 -820
rect 2235 -850 2237 -843
rect 2230 -854 2237 -850
rect 2231 -865 2233 -854
rect 2243 -862 2245 -843
rect 2273 -851 2275 -843
rect 2317 -851 2319 -843
rect 2267 -853 2275 -851
rect 2311 -853 2319 -851
rect 2267 -865 2269 -853
rect 2275 -865 2277 -856
rect 2311 -865 2313 -853
rect 2319 -865 2321 -856
rect 2362 -865 2364 -843
rect 2402 -861 2404 -843
rect 2402 -875 2404 -871
rect 2231 -878 2233 -875
rect 2267 -878 2269 -875
rect 2275 -878 2277 -875
rect 2311 -878 2313 -875
rect 2319 -878 2321 -875
rect 2362 -878 2364 -875
rect 952 -891 956 -890
rect 928 -893 931 -891
rect 941 -893 956 -891
rect 952 -895 956 -893
rect 1059 -891 1063 -890
rect 1035 -893 1038 -891
rect 1048 -893 1063 -891
rect 952 -897 963 -895
rect 988 -897 991 -895
rect 1059 -895 1063 -893
rect 1161 -891 1165 -890
rect 1137 -893 1140 -891
rect 1150 -893 1165 -891
rect 1059 -897 1070 -895
rect 1095 -897 1098 -895
rect 1161 -895 1165 -893
rect 1362 -890 1366 -889
rect 1258 -891 1262 -890
rect 1234 -893 1237 -891
rect 1247 -893 1262 -891
rect 1161 -897 1172 -895
rect 1197 -897 1200 -895
rect 1258 -895 1262 -893
rect 1338 -892 1341 -890
rect 1351 -892 1366 -890
rect 1258 -897 1269 -895
rect 1294 -897 1297 -895
rect 1362 -894 1366 -892
rect 1464 -890 1468 -889
rect 1440 -892 1443 -890
rect 1453 -892 1468 -890
rect 1362 -896 1373 -894
rect 1398 -896 1401 -894
rect 1464 -894 1468 -892
rect 1560 -890 1564 -889
rect 1536 -892 1539 -890
rect 1549 -892 1564 -890
rect 1464 -896 1475 -894
rect 1500 -896 1503 -894
rect 1560 -894 1564 -892
rect 1659 -890 1663 -889
rect 1635 -892 1638 -890
rect 1648 -892 1663 -890
rect 1560 -896 1571 -894
rect 1596 -896 1599 -894
rect 1659 -894 1663 -892
rect 1659 -896 1670 -894
rect 1695 -896 1698 -894
rect 944 -905 963 -903
rect 988 -905 991 -903
rect 1051 -905 1070 -903
rect 1095 -905 1098 -903
rect 1153 -905 1172 -903
rect 1197 -905 1200 -903
rect 1250 -905 1269 -903
rect 1294 -905 1297 -903
rect 1354 -904 1373 -902
rect 1398 -904 1401 -902
rect 1456 -904 1475 -902
rect 1500 -904 1503 -902
rect 1552 -904 1571 -902
rect 1596 -904 1599 -902
rect 1651 -904 1670 -902
rect 1695 -904 1698 -902
rect 928 -929 931 -927
rect 941 -929 955 -927
rect 953 -933 955 -929
rect 1035 -929 1038 -927
rect 1048 -929 1062 -927
rect 953 -935 963 -933
rect 988 -935 991 -933
rect 1060 -933 1062 -929
rect 1137 -929 1140 -927
rect 1150 -929 1164 -927
rect 1060 -935 1070 -933
rect 1095 -935 1098 -933
rect 1162 -933 1164 -929
rect 1234 -929 1237 -927
rect 1247 -929 1261 -927
rect 1338 -928 1341 -926
rect 1351 -928 1365 -926
rect 1162 -935 1172 -933
rect 1197 -935 1200 -933
rect 1259 -933 1261 -929
rect 1259 -935 1269 -933
rect 1294 -935 1297 -933
rect 1363 -932 1365 -928
rect 1440 -928 1443 -926
rect 1453 -928 1467 -926
rect 1363 -934 1373 -932
rect 1398 -934 1401 -932
rect 1465 -932 1467 -928
rect 1536 -928 1539 -926
rect 1549 -928 1563 -926
rect 1465 -934 1475 -932
rect 1500 -934 1503 -932
rect 1561 -932 1563 -928
rect 1635 -928 1638 -926
rect 1648 -928 1662 -926
rect 1561 -934 1571 -932
rect 1596 -934 1599 -932
rect 1660 -932 1662 -928
rect 1660 -934 1670 -932
rect 1695 -934 1698 -932
rect 928 -937 931 -935
rect 941 -937 950 -935
rect 1035 -937 1038 -935
rect 1048 -937 1057 -935
rect 1137 -937 1140 -935
rect 1150 -937 1159 -935
rect 1234 -937 1237 -935
rect 1247 -937 1256 -935
rect 1338 -936 1341 -934
rect 1351 -936 1360 -934
rect 1440 -936 1443 -934
rect 1453 -936 1462 -934
rect 1536 -936 1539 -934
rect 1549 -936 1558 -934
rect 1635 -936 1638 -934
rect 1648 -936 1657 -934
rect 2388 -947 2390 -944
rect 2396 -947 2398 -944
rect 2426 -947 2428 -944
rect 2470 -947 2472 -944
rect 2515 -947 2517 -944
rect 2090 -953 2093 -951
rect 2117 -953 2139 -951
rect 2143 -953 2152 -951
rect 2164 -953 2167 -951
rect 2090 -963 2093 -961
rect 2117 -963 2128 -961
rect 2132 -963 2152 -961
rect 2164 -963 2167 -961
rect 928 -973 931 -971
rect 941 -973 955 -971
rect 953 -977 955 -973
rect 1035 -973 1038 -971
rect 1048 -973 1062 -971
rect 953 -979 963 -977
rect 988 -979 991 -977
rect 1060 -977 1062 -973
rect 1137 -973 1140 -971
rect 1150 -973 1164 -971
rect 1060 -979 1070 -977
rect 1095 -979 1098 -977
rect 1162 -977 1164 -973
rect 1234 -973 1237 -971
rect 1247 -973 1261 -971
rect 1338 -972 1341 -970
rect 1351 -972 1365 -970
rect 1162 -979 1172 -977
rect 1197 -979 1200 -977
rect 1259 -977 1261 -973
rect 1259 -979 1269 -977
rect 1294 -979 1297 -977
rect 1363 -976 1365 -972
rect 1440 -972 1443 -970
rect 1453 -972 1467 -970
rect 1363 -978 1373 -976
rect 1398 -978 1401 -976
rect 1465 -976 1467 -972
rect 1536 -972 1539 -970
rect 1549 -972 1563 -970
rect 1465 -978 1475 -976
rect 1500 -978 1503 -976
rect 1561 -976 1563 -972
rect 1635 -972 1638 -970
rect 1648 -972 1662 -970
rect 1561 -978 1571 -976
rect 1596 -978 1599 -976
rect 1660 -976 1662 -972
rect 2563 -952 2565 -949
rect 1660 -978 1670 -976
rect 1695 -978 1698 -976
rect 928 -981 931 -979
rect 941 -981 950 -979
rect 1035 -981 1038 -979
rect 1048 -981 1057 -979
rect 1137 -981 1140 -979
rect 1150 -981 1159 -979
rect 1234 -981 1237 -979
rect 1247 -981 1256 -979
rect 1338 -980 1341 -978
rect 1351 -980 1360 -978
rect 1440 -980 1443 -978
rect 1453 -980 1462 -978
rect 1536 -980 1539 -978
rect 1549 -980 1558 -978
rect 1635 -980 1638 -978
rect 1648 -980 1657 -978
rect 2388 -979 2390 -972
rect 2084 -981 2087 -979
rect 2111 -981 2121 -979
rect 2126 -981 2152 -979
rect 2164 -981 2167 -979
rect 2084 -991 2087 -989
rect 2111 -991 2120 -989
rect 2383 -983 2390 -979
rect 2125 -991 2152 -989
rect 2164 -991 2167 -989
rect 2384 -994 2386 -983
rect 2396 -991 2398 -972
rect 2426 -980 2428 -972
rect 2470 -980 2472 -972
rect 2420 -982 2428 -980
rect 2464 -982 2472 -980
rect 2420 -994 2422 -982
rect 2428 -994 2430 -985
rect 2464 -994 2466 -982
rect 2472 -994 2474 -985
rect 2515 -994 2517 -972
rect 2563 -990 2565 -972
rect 2259 -1001 2262 -999
rect 2286 -1001 2308 -999
rect 2312 -1001 2321 -999
rect 2333 -1001 2336 -999
rect 2563 -1004 2565 -1000
rect 2384 -1007 2386 -1004
rect 2420 -1007 2422 -1004
rect 2428 -1007 2430 -1004
rect 2464 -1007 2466 -1004
rect 2472 -1007 2474 -1004
rect 2515 -1007 2517 -1004
rect 2259 -1011 2262 -1009
rect 2286 -1011 2297 -1009
rect 2301 -1011 2321 -1009
rect 2333 -1011 2336 -1009
rect 928 -1024 931 -1022
rect 941 -1024 963 -1022
rect 988 -1024 991 -1022
rect 1035 -1024 1038 -1022
rect 1048 -1024 1070 -1022
rect 1095 -1024 1098 -1022
rect 1137 -1024 1140 -1022
rect 1150 -1024 1172 -1022
rect 1197 -1024 1200 -1022
rect 1234 -1024 1237 -1022
rect 1247 -1024 1269 -1022
rect 1294 -1024 1297 -1022
rect 1338 -1023 1341 -1021
rect 1351 -1023 1373 -1021
rect 1398 -1023 1401 -1021
rect 1440 -1023 1443 -1021
rect 1453 -1023 1475 -1021
rect 1500 -1023 1503 -1021
rect 1536 -1023 1539 -1021
rect 1549 -1023 1571 -1021
rect 1596 -1023 1599 -1021
rect 1635 -1023 1638 -1021
rect 1648 -1023 1670 -1021
rect 1695 -1023 1698 -1021
rect 2080 -1030 2083 -1028
rect 2095 -1030 2109 -1028
rect 2115 -1030 2118 -1028
rect 2135 -1030 2138 -1028
rect 2150 -1030 2164 -1028
rect 2170 -1030 2173 -1028
rect 2253 -1029 2256 -1027
rect 2280 -1029 2290 -1027
rect 2295 -1029 2321 -1027
rect 2333 -1029 2336 -1027
rect 2253 -1039 2256 -1037
rect 2280 -1039 2289 -1037
rect 2294 -1039 2321 -1037
rect 2333 -1039 2336 -1037
rect 1716 -1075 1718 -1072
rect 1755 -1079 1757 -1076
rect 1765 -1079 1767 -1076
rect 2249 -1078 2252 -1076
rect 2264 -1078 2278 -1076
rect 2284 -1078 2287 -1076
rect 2304 -1078 2307 -1076
rect 2319 -1078 2333 -1076
rect 2339 -1078 2342 -1076
rect 1716 -1101 1718 -1087
rect 1783 -1085 1785 -1082
rect 1793 -1085 1795 -1082
rect 1716 -1110 1718 -1107
rect 1755 -1112 1757 -1103
rect 1765 -1113 1767 -1103
rect 2582 -1105 2584 -1102
rect 2590 -1105 2592 -1102
rect 2620 -1105 2622 -1102
rect 2664 -1105 2666 -1102
rect 2709 -1105 2711 -1102
rect 1716 -1130 1718 -1127
rect 1716 -1156 1718 -1142
rect 1755 -1144 1757 -1117
rect 1765 -1144 1767 -1118
rect 1783 -1120 1785 -1109
rect 1783 -1144 1785 -1124
rect 1793 -1131 1795 -1109
rect 2756 -1110 2758 -1107
rect 1793 -1144 1795 -1135
rect 2582 -1137 2584 -1130
rect 2577 -1141 2584 -1137
rect 2578 -1152 2580 -1141
rect 2590 -1149 2592 -1130
rect 2620 -1138 2622 -1130
rect 2664 -1138 2666 -1130
rect 2614 -1140 2622 -1138
rect 2658 -1140 2666 -1138
rect 2614 -1152 2616 -1140
rect 2622 -1152 2624 -1143
rect 2658 -1152 2660 -1140
rect 2666 -1152 2668 -1143
rect 2709 -1152 2711 -1130
rect 2756 -1148 2758 -1130
rect 1755 -1159 1757 -1156
rect 1765 -1159 1767 -1156
rect 1783 -1159 1785 -1156
rect 1793 -1159 1795 -1156
rect 2442 -1159 2445 -1157
rect 2469 -1159 2491 -1157
rect 2495 -1159 2504 -1157
rect 2516 -1159 2519 -1157
rect 1716 -1165 1718 -1162
rect 2756 -1162 2758 -1158
rect 2578 -1165 2580 -1162
rect 2614 -1165 2616 -1162
rect 2622 -1165 2624 -1162
rect 2658 -1165 2660 -1162
rect 2666 -1165 2668 -1162
rect 2709 -1165 2711 -1162
rect 2442 -1169 2445 -1167
rect 2469 -1169 2480 -1167
rect 2484 -1169 2504 -1167
rect 2516 -1169 2519 -1167
rect 2436 -1187 2439 -1185
rect 2463 -1187 2473 -1185
rect 2478 -1187 2504 -1185
rect 2516 -1187 2519 -1185
rect 2436 -1197 2439 -1195
rect 2463 -1197 2472 -1195
rect 2477 -1197 2504 -1195
rect 2516 -1197 2519 -1195
rect 1717 -1207 1719 -1204
rect 1756 -1211 1758 -1208
rect 1766 -1211 1768 -1208
rect 1717 -1233 1719 -1219
rect 1784 -1217 1786 -1214
rect 1794 -1217 1796 -1214
rect 1717 -1242 1719 -1239
rect 1756 -1244 1758 -1235
rect 1766 -1245 1768 -1235
rect 2432 -1236 2435 -1234
rect 2447 -1236 2461 -1234
rect 2467 -1236 2470 -1234
rect 2487 -1236 2490 -1234
rect 2502 -1236 2516 -1234
rect 2522 -1236 2525 -1234
rect 1717 -1262 1719 -1259
rect 1717 -1288 1719 -1274
rect 1756 -1276 1758 -1249
rect 1766 -1276 1768 -1250
rect 1784 -1252 1786 -1241
rect 1784 -1276 1786 -1256
rect 1794 -1263 1796 -1241
rect 2053 -1252 2056 -1250
rect 2096 -1252 2114 -1250
rect 2134 -1252 2138 -1250
rect 1794 -1276 1796 -1267
rect 1756 -1291 1758 -1288
rect 1766 -1291 1768 -1288
rect 1784 -1291 1786 -1288
rect 1794 -1291 1796 -1288
rect 1717 -1297 1719 -1294
rect 2220 -1295 2223 -1293
rect 2263 -1295 2281 -1293
rect 2301 -1295 2305 -1293
rect 2402 -1302 2405 -1300
rect 2445 -1302 2463 -1300
rect 2483 -1302 2487 -1300
rect 1720 -1351 1722 -1348
rect 1759 -1355 1761 -1352
rect 1769 -1355 1771 -1352
rect 1720 -1377 1722 -1363
rect 1787 -1361 1789 -1358
rect 1797 -1361 1799 -1358
rect 1720 -1386 1722 -1383
rect 1759 -1388 1761 -1379
rect 1769 -1389 1771 -1379
rect 1720 -1406 1722 -1403
rect 1720 -1432 1722 -1418
rect 1759 -1420 1761 -1393
rect 1769 -1420 1771 -1394
rect 1787 -1396 1789 -1385
rect 1787 -1420 1789 -1400
rect 1797 -1407 1799 -1385
rect 2696 -1391 2698 -1388
rect 1797 -1420 1799 -1411
rect 2743 -1410 2745 -1407
rect 2751 -1410 2753 -1407
rect 2781 -1410 2783 -1407
rect 2825 -1410 2827 -1407
rect 2870 -1410 2872 -1407
rect 1759 -1435 1761 -1432
rect 1769 -1435 1771 -1432
rect 1787 -1435 1789 -1432
rect 1797 -1435 1799 -1432
rect 1720 -1441 1722 -1438
rect 2696 -1449 2698 -1431
rect 2908 -1418 2910 -1415
rect 2743 -1442 2745 -1435
rect 2738 -1446 2745 -1442
rect 2559 -1457 2562 -1455
rect 2612 -1457 2635 -1455
rect 2739 -1457 2741 -1446
rect 2751 -1454 2753 -1435
rect 2781 -1443 2783 -1435
rect 2825 -1443 2827 -1435
rect 2775 -1445 2783 -1443
rect 2819 -1445 2827 -1443
rect 2775 -1457 2777 -1445
rect 2783 -1457 2785 -1448
rect 2819 -1457 2821 -1445
rect 2827 -1457 2829 -1448
rect 2870 -1457 2872 -1435
rect 2908 -1456 2910 -1438
rect 2696 -1473 2698 -1469
rect 2739 -1470 2741 -1467
rect 2775 -1470 2777 -1467
rect 2783 -1470 2785 -1467
rect 2819 -1470 2821 -1467
rect 2827 -1470 2829 -1467
rect 2870 -1470 2872 -1467
rect 2908 -1470 2910 -1466
rect 1727 -1476 1729 -1473
rect 1766 -1480 1768 -1477
rect 1776 -1480 1778 -1477
rect 1727 -1502 1729 -1488
rect 1794 -1486 1796 -1483
rect 1804 -1486 1806 -1483
rect 1727 -1511 1729 -1508
rect 1766 -1513 1768 -1504
rect 1776 -1514 1778 -1504
rect 2363 -1492 2366 -1490
rect 2416 -1492 2439 -1490
rect 2189 -1496 2192 -1494
rect 2242 -1496 2265 -1494
rect 1727 -1531 1729 -1528
rect 1727 -1557 1729 -1543
rect 1766 -1545 1768 -1518
rect 1776 -1545 1778 -1519
rect 1794 -1521 1796 -1510
rect 1794 -1545 1796 -1525
rect 1804 -1532 1806 -1510
rect 2015 -1519 2018 -1517
rect 2068 -1519 2091 -1517
rect 1804 -1545 1806 -1536
rect 2526 -1542 2538 -1540
rect 2638 -1542 2641 -1540
rect 2338 -1550 2350 -1548
rect 2450 -1550 2453 -1548
rect 1766 -1560 1768 -1557
rect 1776 -1560 1778 -1557
rect 1794 -1560 1796 -1557
rect 1804 -1560 1806 -1557
rect 2157 -1560 2169 -1558
rect 2269 -1560 2272 -1558
rect 1727 -1566 1729 -1563
rect 1989 -1568 2001 -1566
rect 2101 -1568 2104 -1566
rect 2528 -1651 2540 -1649
rect 2640 -1651 2643 -1649
rect 2336 -1661 2348 -1659
rect 2448 -1661 2451 -1659
rect 2156 -1671 2168 -1669
rect 2268 -1671 2271 -1669
rect 1953 -1679 1955 -1676
rect 1749 -1701 1751 -1698
rect 1760 -1701 1762 -1698
rect 1791 -1708 1793 -1704
rect 1749 -1750 1751 -1721
rect 1760 -1750 1762 -1721
rect 1791 -1742 1793 -1728
rect 1791 -1755 1793 -1752
rect 1749 -1773 1751 -1770
rect 1760 -1773 1762 -1770
rect 1988 -1682 2000 -1680
rect 2100 -1682 2103 -1680
rect 1953 -1791 1955 -1779
rect 2030 -1780 2033 -1778
rect 2133 -1780 2145 -1778
rect 1749 -1810 1751 -1807
rect 1760 -1810 1762 -1807
rect 2087 -1811 2090 -1809
rect 2130 -1811 2148 -1809
rect 2168 -1811 2172 -1809
rect 1791 -1817 1793 -1813
rect 1749 -1859 1751 -1830
rect 1760 -1859 1762 -1830
rect 1791 -1851 1793 -1837
rect 1896 -1840 1899 -1838
rect 1924 -1840 1946 -1838
rect 1956 -1840 1959 -1838
rect 1791 -1864 1793 -1861
rect 1749 -1882 1751 -1879
rect 1760 -1882 1762 -1879
rect 1937 -1883 1946 -1881
rect 1956 -1883 1959 -1881
rect 1896 -1885 1899 -1883
rect 1924 -1885 1934 -1883
rect 1932 -1889 1934 -1885
rect 1932 -1891 1946 -1889
rect 1956 -1891 1959 -1889
rect 1750 -1929 1752 -1926
rect 1761 -1929 1763 -1926
rect 1937 -1927 1946 -1925
rect 1956 -1927 1959 -1925
rect 1896 -1929 1899 -1927
rect 1924 -1929 1934 -1927
rect 1792 -1936 1794 -1932
rect 1932 -1933 1934 -1929
rect 1932 -1935 1946 -1933
rect 1956 -1935 1959 -1933
rect 1750 -1978 1752 -1949
rect 1761 -1978 1763 -1949
rect 1792 -1970 1794 -1956
rect 1896 -1959 1899 -1957
rect 1924 -1959 1943 -1957
rect 1896 -1967 1899 -1965
rect 1924 -1967 1935 -1965
rect 1931 -1969 1935 -1967
rect 1931 -1971 1946 -1969
rect 1956 -1971 1959 -1969
rect 1931 -1972 1935 -1971
rect 1792 -1983 1794 -1980
rect 1750 -2001 1752 -1998
rect 1761 -2001 1763 -1998
rect 1754 -2037 1756 -2034
rect 1765 -2037 1767 -2034
rect 1796 -2044 1798 -2040
rect 1754 -2086 1756 -2057
rect 1765 -2086 1767 -2057
rect 1796 -2078 1798 -2064
rect 1796 -2091 1798 -2088
rect 1754 -2109 1756 -2106
rect 1765 -2109 1767 -2106
<< polycontact >>
rect 2077 -703 2081 -699
rect 2077 -758 2081 -754
rect 2146 -729 2150 -725
rect 2157 -740 2161 -736
rect 2212 -750 2216 -746
rect 2225 -758 2229 -754
rect 2236 -750 2240 -746
rect 2248 -758 2253 -753
rect 2263 -758 2267 -754
rect 2292 -758 2297 -753
rect 2344 -753 2348 -748
rect 2307 -758 2311 -754
rect 2226 -854 2230 -850
rect 2239 -862 2243 -858
rect 2250 -854 2254 -850
rect 2262 -862 2267 -857
rect 2277 -862 2281 -858
rect 2306 -862 2311 -857
rect 2358 -857 2362 -852
rect 2321 -862 2325 -858
rect 952 -890 956 -886
rect 1059 -890 1063 -886
rect 1161 -890 1165 -886
rect 1258 -890 1262 -886
rect 1362 -889 1366 -885
rect 1464 -889 1468 -885
rect 1560 -889 1564 -885
rect 1659 -889 1663 -885
rect 944 -903 948 -899
rect 1051 -903 1055 -899
rect 1153 -903 1157 -899
rect 1250 -903 1254 -899
rect 1354 -902 1358 -898
rect 1456 -902 1460 -898
rect 1552 -902 1556 -898
rect 1651 -902 1655 -898
rect 952 -914 956 -910
rect 1059 -914 1063 -910
rect 1161 -914 1165 -910
rect 1258 -914 1262 -910
rect 1362 -913 1366 -909
rect 1464 -913 1468 -909
rect 1560 -913 1564 -909
rect 1659 -913 1663 -909
rect 944 -927 949 -922
rect 1051 -927 1056 -922
rect 1153 -927 1158 -922
rect 1250 -927 1255 -922
rect 1354 -926 1359 -921
rect 1456 -926 1461 -921
rect 1552 -926 1557 -921
rect 1651 -926 1656 -921
rect 944 -941 948 -937
rect 1051 -941 1055 -937
rect 1153 -941 1157 -937
rect 1250 -941 1254 -937
rect 1354 -940 1358 -936
rect 1456 -940 1460 -936
rect 1552 -940 1556 -936
rect 1651 -940 1655 -936
rect 2139 -954 2143 -950
rect 944 -971 949 -966
rect 1051 -971 1056 -966
rect 1153 -971 1158 -966
rect 1250 -971 1255 -966
rect 1354 -970 1359 -965
rect 1456 -970 1461 -965
rect 1552 -970 1557 -965
rect 1651 -970 1656 -965
rect 2128 -965 2132 -961
rect 944 -985 948 -981
rect 1051 -985 1055 -981
rect 1153 -985 1157 -981
rect 1250 -985 1254 -981
rect 1354 -984 1358 -980
rect 1456 -984 1460 -980
rect 1552 -984 1556 -980
rect 1651 -984 1655 -980
rect 2379 -983 2383 -979
rect 2392 -991 2396 -987
rect 2403 -983 2407 -979
rect 2415 -991 2420 -986
rect 2430 -991 2434 -987
rect 2459 -991 2464 -986
rect 2511 -986 2515 -981
rect 2474 -991 2478 -987
rect 2308 -1002 2312 -998
rect 2297 -1013 2301 -1009
rect 949 -1022 954 -1018
rect 1056 -1022 1061 -1018
rect 1158 -1022 1163 -1018
rect 1255 -1022 1260 -1018
rect 1359 -1021 1364 -1017
rect 1461 -1021 1466 -1017
rect 1557 -1021 1562 -1017
rect 1656 -1021 1661 -1017
rect 2102 -1034 2106 -1030
rect 2157 -1034 2161 -1030
rect 1712 -1098 1716 -1094
rect 2271 -1082 2275 -1078
rect 2326 -1082 2330 -1078
rect 1712 -1153 1716 -1149
rect 1781 -1124 1785 -1120
rect 1792 -1135 1796 -1131
rect 2573 -1141 2577 -1137
rect 2586 -1149 2590 -1145
rect 2597 -1141 2601 -1137
rect 2609 -1149 2614 -1144
rect 2624 -1149 2628 -1145
rect 2653 -1149 2658 -1144
rect 2705 -1144 2709 -1139
rect 2668 -1149 2672 -1145
rect 2491 -1160 2495 -1156
rect 2480 -1171 2484 -1167
rect 1713 -1230 1717 -1226
rect 2454 -1240 2458 -1236
rect 2509 -1240 2513 -1236
rect 1713 -1285 1717 -1281
rect 1782 -1256 1786 -1252
rect 1793 -1267 1797 -1263
rect 1716 -1374 1720 -1370
rect 1716 -1429 1720 -1425
rect 1785 -1400 1789 -1396
rect 1796 -1411 1800 -1407
rect 2691 -1446 2696 -1441
rect 2734 -1446 2738 -1442
rect 2747 -1454 2751 -1450
rect 2758 -1446 2762 -1442
rect 2770 -1454 2775 -1449
rect 2785 -1454 2789 -1450
rect 2814 -1454 2819 -1449
rect 2866 -1449 2870 -1444
rect 2829 -1454 2833 -1450
rect 1723 -1499 1727 -1495
rect 1723 -1554 1727 -1550
rect 1792 -1525 1796 -1521
rect 1803 -1536 1807 -1532
rect 1745 -1747 1749 -1743
rect 1756 -1740 1760 -1736
rect 1787 -1739 1791 -1735
rect 1745 -1856 1749 -1852
rect 1756 -1849 1760 -1845
rect 1787 -1848 1791 -1844
rect 1933 -1844 1938 -1840
rect 1939 -1881 1943 -1877
rect 1938 -1896 1943 -1891
rect 1939 -1925 1943 -1921
rect 1746 -1975 1750 -1971
rect 1757 -1968 1761 -1964
rect 1938 -1940 1943 -1935
rect 1931 -1952 1935 -1948
rect 1788 -1967 1792 -1963
rect 1939 -1963 1943 -1959
rect 1931 -1976 1935 -1972
rect 1750 -2083 1754 -2079
rect 1761 -2076 1765 -2072
rect 1792 -2075 1796 -2071
<< metal1 >>
rect 2075 -674 2103 -671
rect 2076 -680 2079 -674
rect 2100 -675 2103 -674
rect 2100 -678 2171 -675
rect 1915 -704 2062 -701
rect 922 -886 926 -885
rect 922 -890 931 -886
rect 952 -886 956 -879
rect 994 -890 998 -884
rect 922 -922 926 -890
rect 931 -906 941 -898
rect 944 -899 948 -890
rect 988 -894 998 -890
rect 931 -910 963 -906
rect 947 -919 949 -914
rect 944 -922 949 -919
rect 952 -915 956 -914
rect 922 -926 931 -922
rect 922 -966 926 -926
rect 994 -928 998 -894
rect 988 -932 998 -928
rect 931 -950 941 -942
rect 944 -942 948 -941
rect 963 -950 988 -940
rect 931 -953 988 -950
rect 949 -958 954 -953
rect 944 -962 954 -958
rect 944 -966 949 -962
rect 922 -970 931 -966
rect 922 -1017 926 -970
rect 994 -972 998 -932
rect 988 -976 998 -972
rect 931 -994 941 -986
rect 944 -986 948 -985
rect 963 -994 988 -984
rect 931 -997 988 -994
rect 922 -1021 931 -1017
rect 949 -1018 954 -997
rect 994 -1017 998 -976
rect 922 -1029 926 -1021
rect 988 -1021 998 -1017
rect 941 -1029 963 -1025
rect 948 -1032 953 -1029
rect 994 -1037 998 -1021
rect 1029 -886 1033 -885
rect 1029 -890 1038 -886
rect 1059 -886 1063 -879
rect 1101 -890 1105 -884
rect 1029 -922 1033 -890
rect 1038 -906 1048 -898
rect 1051 -899 1055 -890
rect 1095 -894 1105 -890
rect 1038 -910 1070 -906
rect 1054 -919 1056 -914
rect 1051 -922 1056 -919
rect 1059 -915 1063 -914
rect 1029 -926 1038 -922
rect 1029 -966 1033 -926
rect 1101 -928 1105 -894
rect 1095 -932 1105 -928
rect 1038 -950 1048 -942
rect 1051 -942 1055 -941
rect 1070 -950 1095 -940
rect 1038 -953 1095 -950
rect 1056 -958 1061 -953
rect 1051 -962 1061 -958
rect 1051 -966 1056 -962
rect 1029 -970 1038 -966
rect 1029 -1017 1033 -970
rect 1101 -972 1105 -932
rect 1095 -976 1105 -972
rect 1038 -994 1048 -986
rect 1051 -986 1055 -985
rect 1070 -994 1095 -984
rect 1038 -997 1095 -994
rect 1029 -1021 1038 -1017
rect 1056 -1018 1061 -997
rect 1101 -1017 1105 -976
rect 1029 -1029 1033 -1021
rect 1095 -1021 1105 -1017
rect 1048 -1029 1070 -1025
rect 1055 -1032 1060 -1029
rect 1101 -1037 1105 -1021
rect 1131 -886 1135 -885
rect 1131 -890 1140 -886
rect 1161 -886 1165 -879
rect 1203 -890 1207 -884
rect 1131 -922 1135 -890
rect 1140 -906 1150 -898
rect 1153 -899 1157 -890
rect 1197 -894 1207 -890
rect 1140 -910 1172 -906
rect 1156 -919 1158 -914
rect 1153 -922 1158 -919
rect 1161 -915 1165 -914
rect 1131 -926 1140 -922
rect 1131 -966 1135 -926
rect 1203 -928 1207 -894
rect 1197 -932 1207 -928
rect 1140 -950 1150 -942
rect 1153 -942 1157 -941
rect 1172 -950 1197 -940
rect 1140 -953 1197 -950
rect 1158 -958 1163 -953
rect 1153 -962 1163 -958
rect 1153 -966 1158 -962
rect 1131 -970 1140 -966
rect 1131 -1017 1135 -970
rect 1203 -972 1207 -932
rect 1197 -976 1207 -972
rect 1140 -994 1150 -986
rect 1153 -986 1157 -985
rect 1172 -994 1197 -984
rect 1140 -997 1197 -994
rect 1131 -1021 1140 -1017
rect 1158 -1018 1163 -997
rect 1203 -1017 1207 -976
rect 1131 -1029 1135 -1021
rect 1197 -1021 1207 -1017
rect 1150 -1029 1172 -1025
rect 1157 -1032 1162 -1029
rect 1203 -1037 1207 -1021
rect 1228 -886 1232 -885
rect 1228 -890 1237 -886
rect 1258 -886 1262 -879
rect 1300 -890 1304 -884
rect 1228 -922 1232 -890
rect 1237 -906 1247 -898
rect 1250 -899 1254 -890
rect 1294 -894 1304 -890
rect 1237 -910 1269 -906
rect 1253 -919 1255 -914
rect 1250 -922 1255 -919
rect 1258 -915 1262 -914
rect 1228 -926 1237 -922
rect 1228 -966 1232 -926
rect 1300 -928 1304 -894
rect 1294 -932 1304 -928
rect 1237 -950 1247 -942
rect 1250 -942 1254 -941
rect 1269 -950 1294 -940
rect 1237 -953 1294 -950
rect 1255 -958 1260 -953
rect 1250 -962 1260 -958
rect 1250 -966 1255 -962
rect 1228 -970 1237 -966
rect 1228 -1017 1232 -970
rect 1300 -972 1304 -932
rect 1294 -976 1304 -972
rect 1237 -994 1247 -986
rect 1250 -986 1254 -985
rect 1269 -994 1294 -984
rect 1237 -997 1294 -994
rect 1228 -1021 1237 -1017
rect 1255 -1018 1260 -997
rect 1300 -1017 1304 -976
rect 1228 -1029 1232 -1021
rect 1294 -1021 1304 -1017
rect 1247 -1029 1269 -1025
rect 1254 -1032 1259 -1029
rect 1300 -1037 1304 -1021
rect 1332 -885 1336 -884
rect 1332 -889 1341 -885
rect 1362 -885 1366 -878
rect 1404 -889 1408 -883
rect 1332 -921 1336 -889
rect 1341 -905 1351 -897
rect 1354 -898 1358 -889
rect 1398 -893 1408 -889
rect 1341 -909 1373 -905
rect 1357 -918 1359 -913
rect 1354 -921 1359 -918
rect 1362 -914 1366 -913
rect 1332 -925 1341 -921
rect 1332 -965 1336 -925
rect 1404 -927 1408 -893
rect 1398 -931 1408 -927
rect 1341 -949 1351 -941
rect 1354 -941 1358 -940
rect 1373 -949 1398 -939
rect 1341 -952 1398 -949
rect 1359 -957 1364 -952
rect 1354 -961 1364 -957
rect 1354 -965 1359 -961
rect 1332 -969 1341 -965
rect 1332 -1016 1336 -969
rect 1404 -971 1408 -931
rect 1398 -975 1408 -971
rect 1341 -993 1351 -985
rect 1354 -985 1358 -984
rect 1373 -993 1398 -983
rect 1341 -996 1398 -993
rect 1332 -1020 1341 -1016
rect 1359 -1017 1364 -996
rect 1404 -1016 1408 -975
rect 1332 -1028 1336 -1020
rect 1398 -1020 1408 -1016
rect 1351 -1028 1373 -1024
rect 1358 -1031 1363 -1028
rect 1404 -1036 1408 -1020
rect 1434 -885 1438 -884
rect 1434 -889 1443 -885
rect 1464 -885 1468 -878
rect 1506 -889 1510 -883
rect 1434 -921 1438 -889
rect 1443 -905 1453 -897
rect 1456 -898 1460 -889
rect 1500 -893 1510 -889
rect 1443 -909 1475 -905
rect 1459 -918 1461 -913
rect 1456 -921 1461 -918
rect 1464 -914 1468 -913
rect 1434 -925 1443 -921
rect 1434 -965 1438 -925
rect 1506 -927 1510 -893
rect 1500 -931 1510 -927
rect 1443 -949 1453 -941
rect 1456 -941 1460 -940
rect 1475 -949 1500 -939
rect 1443 -952 1500 -949
rect 1461 -957 1466 -952
rect 1456 -961 1466 -957
rect 1456 -965 1461 -961
rect 1434 -969 1443 -965
rect 1434 -1016 1438 -969
rect 1506 -971 1510 -931
rect 1500 -975 1510 -971
rect 1443 -993 1453 -985
rect 1456 -985 1460 -984
rect 1475 -993 1500 -983
rect 1443 -996 1500 -993
rect 1434 -1020 1443 -1016
rect 1461 -1017 1466 -996
rect 1506 -1016 1510 -975
rect 1434 -1028 1438 -1020
rect 1500 -1020 1510 -1016
rect 1453 -1028 1475 -1024
rect 1460 -1031 1465 -1028
rect 1506 -1036 1510 -1020
rect 1530 -885 1534 -884
rect 1530 -889 1539 -885
rect 1560 -885 1564 -878
rect 1602 -889 1606 -883
rect 1530 -921 1534 -889
rect 1539 -905 1549 -897
rect 1552 -898 1556 -889
rect 1596 -893 1606 -889
rect 1539 -909 1571 -905
rect 1555 -918 1557 -913
rect 1552 -921 1557 -918
rect 1560 -914 1564 -913
rect 1530 -925 1539 -921
rect 1530 -965 1534 -925
rect 1602 -927 1606 -893
rect 1596 -931 1606 -927
rect 1539 -949 1549 -941
rect 1552 -941 1556 -940
rect 1571 -949 1596 -939
rect 1539 -952 1596 -949
rect 1557 -957 1562 -952
rect 1552 -961 1562 -957
rect 1552 -965 1557 -961
rect 1530 -969 1539 -965
rect 1530 -1016 1534 -969
rect 1602 -971 1606 -931
rect 1596 -975 1606 -971
rect 1539 -993 1549 -985
rect 1552 -985 1556 -984
rect 1571 -993 1596 -983
rect 1539 -996 1596 -993
rect 1530 -1020 1539 -1016
rect 1557 -1017 1562 -996
rect 1602 -1016 1606 -975
rect 1530 -1028 1534 -1020
rect 1596 -1020 1606 -1016
rect 1549 -1028 1571 -1024
rect 1556 -1031 1561 -1028
rect 1602 -1036 1606 -1020
rect 1629 -885 1633 -884
rect 1629 -889 1638 -885
rect 1659 -885 1663 -878
rect 1701 -889 1705 -883
rect 1629 -921 1633 -889
rect 1638 -905 1648 -897
rect 1651 -898 1655 -889
rect 1695 -893 1705 -889
rect 1638 -909 1670 -905
rect 1654 -918 1656 -913
rect 1651 -921 1656 -918
rect 1659 -914 1663 -913
rect 1629 -925 1638 -921
rect 1629 -965 1633 -925
rect 1701 -927 1705 -893
rect 1695 -931 1705 -927
rect 1638 -949 1648 -941
rect 1651 -941 1655 -940
rect 1670 -949 1695 -939
rect 1638 -952 1695 -949
rect 1656 -957 1661 -952
rect 1651 -961 1661 -957
rect 1651 -965 1656 -961
rect 1629 -969 1638 -965
rect 1629 -1016 1633 -969
rect 1701 -971 1705 -931
rect 1695 -975 1705 -971
rect 1638 -993 1648 -985
rect 1651 -985 1655 -984
rect 1670 -993 1695 -983
rect 1638 -996 1695 -993
rect 1629 -1020 1638 -1016
rect 1656 -1017 1661 -996
rect 1701 -1016 1705 -975
rect 1629 -1028 1633 -1020
rect 1695 -1020 1705 -1016
rect 1648 -1028 1670 -1024
rect 1655 -1030 1660 -1028
rect 1701 -1036 1705 -1020
rect 1655 -1037 1660 -1036
rect 1710 -1069 1738 -1066
rect 1711 -1075 1714 -1069
rect 1735 -1070 1738 -1069
rect 1735 -1073 1806 -1070
rect 948 -1099 1655 -1096
rect 1660 -1099 1697 -1096
rect 1702 -1098 1712 -1095
rect 1720 -1095 1723 -1087
rect 1750 -1079 1753 -1073
rect 1769 -1079 1772 -1073
rect 1720 -1098 1741 -1095
rect 1720 -1101 1723 -1098
rect 1711 -1111 1714 -1107
rect 1705 -1113 1729 -1111
rect 1705 -1114 1723 -1113
rect 1728 -1114 1729 -1113
rect 1738 -1121 1741 -1098
rect 1779 -1079 1799 -1076
rect 1779 -1085 1782 -1079
rect 1796 -1085 1799 -1079
rect 1760 -1106 1763 -1103
rect 1760 -1109 1778 -1106
rect 1788 -1116 1791 -1109
rect 1788 -1119 1805 -1116
rect 1710 -1122 1729 -1121
rect 1705 -1124 1729 -1122
rect 1738 -1124 1781 -1121
rect 1711 -1130 1714 -1124
rect 1802 -1130 1805 -1119
rect 1767 -1135 1792 -1132
rect 1802 -1134 1815 -1130
rect 1767 -1137 1770 -1135
rect 948 -1153 1556 -1150
rect 1561 -1153 1697 -1150
rect 1702 -1153 1712 -1150
rect 1720 -1150 1723 -1142
rect 1732 -1140 1770 -1137
rect 1802 -1138 1805 -1134
rect 1732 -1150 1735 -1140
rect 1773 -1141 1805 -1138
rect 1773 -1144 1776 -1141
rect 1720 -1153 1735 -1150
rect 1720 -1156 1723 -1153
rect 1772 -1147 1778 -1144
rect 1711 -1166 1714 -1162
rect 1732 -1163 1737 -1160
rect 1750 -1160 1753 -1156
rect 1797 -1160 1800 -1156
rect 1742 -1163 1806 -1160
rect 1732 -1166 1735 -1163
rect 1705 -1169 1735 -1166
rect 1811 -1169 1815 -1134
rect 1711 -1201 1739 -1198
rect 1712 -1207 1715 -1201
rect 1736 -1202 1739 -1201
rect 1736 -1205 1807 -1202
rect 948 -1231 1460 -1228
rect 1465 -1231 1698 -1228
rect 1703 -1230 1713 -1227
rect 1721 -1227 1724 -1219
rect 1751 -1211 1754 -1205
rect 1770 -1211 1773 -1205
rect 1721 -1230 1742 -1227
rect 1721 -1233 1724 -1230
rect 1712 -1243 1715 -1239
rect 1706 -1245 1730 -1243
rect 1706 -1246 1724 -1245
rect 1729 -1246 1730 -1245
rect 1739 -1253 1742 -1230
rect 1780 -1211 1800 -1208
rect 1780 -1217 1783 -1211
rect 1797 -1217 1800 -1211
rect 1761 -1238 1764 -1235
rect 1761 -1241 1779 -1238
rect 1789 -1248 1792 -1241
rect 1789 -1251 1806 -1248
rect 1711 -1254 1730 -1253
rect 1706 -1256 1730 -1254
rect 1739 -1256 1782 -1253
rect 1712 -1262 1715 -1256
rect 1803 -1262 1806 -1251
rect 1768 -1267 1793 -1264
rect 1803 -1266 1816 -1262
rect 1768 -1269 1771 -1267
rect 948 -1285 1358 -1282
rect 1363 -1285 1698 -1282
rect 1703 -1285 1713 -1282
rect 1721 -1282 1724 -1274
rect 1733 -1272 1771 -1269
rect 1803 -1270 1806 -1266
rect 1733 -1282 1736 -1272
rect 1774 -1273 1806 -1270
rect 1774 -1276 1777 -1273
rect 1721 -1285 1736 -1282
rect 1721 -1288 1724 -1285
rect 1773 -1279 1779 -1276
rect 1712 -1298 1715 -1294
rect 1733 -1295 1738 -1292
rect 1751 -1292 1754 -1288
rect 1798 -1292 1801 -1288
rect 1743 -1295 1807 -1292
rect 1733 -1298 1736 -1295
rect 1706 -1301 1736 -1298
rect 1812 -1299 1816 -1266
rect 1812 -1306 1816 -1304
rect 1714 -1345 1742 -1342
rect 1715 -1351 1718 -1345
rect 1739 -1346 1742 -1345
rect 1739 -1349 1810 -1346
rect 948 -1375 1254 -1372
rect 1259 -1375 1701 -1372
rect 1706 -1374 1716 -1371
rect 1724 -1371 1727 -1363
rect 1754 -1355 1757 -1349
rect 1773 -1355 1776 -1349
rect 1724 -1374 1745 -1371
rect 1724 -1377 1727 -1374
rect 1715 -1387 1718 -1383
rect 1709 -1389 1733 -1387
rect 1709 -1390 1727 -1389
rect 1732 -1390 1733 -1389
rect 1742 -1397 1745 -1374
rect 1783 -1355 1803 -1352
rect 1783 -1361 1786 -1355
rect 1800 -1361 1803 -1355
rect 1764 -1382 1767 -1379
rect 1764 -1385 1782 -1382
rect 1792 -1392 1795 -1385
rect 1792 -1395 1809 -1392
rect 1714 -1398 1733 -1397
rect 1709 -1400 1733 -1398
rect 1742 -1400 1785 -1397
rect 1715 -1406 1718 -1400
rect 1806 -1406 1809 -1395
rect 1771 -1411 1796 -1408
rect 1806 -1410 1819 -1406
rect 1771 -1413 1774 -1411
rect 948 -1429 1157 -1426
rect 1162 -1429 1701 -1426
rect 1706 -1429 1716 -1426
rect 1724 -1426 1727 -1418
rect 1736 -1416 1774 -1413
rect 1806 -1414 1809 -1410
rect 1736 -1426 1739 -1416
rect 1777 -1417 1809 -1414
rect 1777 -1420 1780 -1417
rect 1724 -1429 1739 -1426
rect 1724 -1432 1727 -1429
rect 1776 -1423 1782 -1420
rect 1715 -1442 1718 -1438
rect 1736 -1439 1741 -1436
rect 1754 -1436 1757 -1432
rect 1801 -1436 1804 -1432
rect 1746 -1439 1810 -1436
rect 1736 -1442 1739 -1439
rect 1709 -1445 1739 -1442
rect 1815 -1445 1819 -1410
rect 1721 -1470 1749 -1467
rect 1722 -1476 1725 -1470
rect 1746 -1471 1749 -1470
rect 1746 -1474 1817 -1471
rect 948 -1500 1055 -1497
rect 1060 -1500 1708 -1497
rect 1713 -1499 1723 -1496
rect 1731 -1496 1734 -1488
rect 1761 -1480 1764 -1474
rect 1780 -1480 1783 -1474
rect 1731 -1499 1752 -1496
rect 1731 -1502 1734 -1499
rect 1722 -1512 1725 -1508
rect 1716 -1514 1740 -1512
rect 1716 -1515 1734 -1514
rect 1739 -1515 1740 -1514
rect 1749 -1522 1752 -1499
rect 1790 -1480 1810 -1477
rect 1790 -1486 1793 -1480
rect 1807 -1486 1810 -1480
rect 1771 -1507 1774 -1504
rect 1771 -1510 1789 -1507
rect 1799 -1517 1802 -1510
rect 1799 -1520 1816 -1517
rect 1721 -1523 1740 -1522
rect 1716 -1525 1740 -1523
rect 1749 -1525 1792 -1522
rect 1722 -1531 1725 -1525
rect 1813 -1531 1816 -1520
rect 1778 -1536 1803 -1533
rect 1813 -1535 1826 -1531
rect 1778 -1538 1781 -1536
rect 953 -1554 1708 -1551
rect 1713 -1554 1723 -1551
rect 1731 -1551 1734 -1543
rect 1743 -1541 1781 -1538
rect 1813 -1539 1816 -1535
rect 1743 -1551 1746 -1541
rect 1784 -1542 1816 -1539
rect 1784 -1545 1787 -1542
rect 1731 -1554 1746 -1551
rect 1731 -1557 1734 -1554
rect 1783 -1548 1789 -1545
rect 1722 -1567 1725 -1563
rect 1743 -1564 1748 -1561
rect 1761 -1561 1764 -1557
rect 1808 -1561 1811 -1557
rect 1753 -1564 1817 -1561
rect 1743 -1567 1746 -1564
rect 1716 -1570 1746 -1567
rect 1822 -1572 1826 -1535
rect 1744 -1690 1767 -1686
rect 1748 -1692 1767 -1690
rect 1744 -1701 1748 -1696
rect 1763 -1701 1767 -1692
rect 1780 -1697 1804 -1696
rect 1780 -1701 1796 -1697
rect 1800 -1701 1804 -1697
rect 1780 -1703 1804 -1701
rect 1786 -1708 1790 -1703
rect 1755 -1729 1759 -1721
rect 1755 -1733 1767 -1729
rect 1763 -1735 1767 -1733
rect 1794 -1735 1798 -1728
rect 948 -1740 1055 -1736
rect 1060 -1740 1756 -1736
rect 1763 -1739 1787 -1735
rect 1794 -1739 1817 -1735
rect 953 -1747 1745 -1743
rect 1763 -1750 1767 -1739
rect 1794 -1742 1798 -1739
rect 1801 -1740 1817 -1739
rect 1786 -1756 1790 -1752
rect 1780 -1757 1805 -1756
rect 1780 -1761 1800 -1757
rect 1780 -1762 1805 -1761
rect 1744 -1774 1748 -1770
rect 1744 -1778 1760 -1774
rect 1915 -1778 1918 -704
rect 2067 -703 2077 -700
rect 2085 -700 2088 -692
rect 2115 -684 2118 -678
rect 2134 -684 2137 -678
rect 2085 -703 2106 -700
rect 2085 -706 2088 -703
rect 2076 -716 2079 -712
rect 2070 -718 2094 -716
rect 2070 -719 2088 -718
rect 2093 -719 2094 -718
rect 2103 -726 2106 -703
rect 2144 -684 2164 -681
rect 2144 -690 2147 -684
rect 2161 -690 2164 -684
rect 2125 -711 2128 -708
rect 2125 -714 2143 -711
rect 2210 -708 2363 -704
rect 2216 -714 2220 -708
rect 2254 -714 2258 -708
rect 2298 -714 2302 -708
rect 2343 -714 2347 -708
rect 2392 -709 2396 -706
rect 2386 -713 2387 -709
rect 2391 -713 2396 -709
rect 2153 -721 2156 -714
rect 2153 -724 2170 -721
rect 2075 -727 2094 -726
rect 2070 -729 2094 -727
rect 2103 -729 2146 -726
rect 2076 -735 2079 -729
rect 2167 -735 2170 -724
rect 2132 -740 2157 -737
rect 2167 -739 2180 -735
rect 2266 -739 2279 -714
rect 2310 -739 2323 -714
rect 2392 -719 2396 -713
rect 2132 -742 2135 -740
rect 1994 -758 2062 -753
rect 2067 -758 2077 -755
rect 2085 -755 2088 -747
rect 2097 -745 2135 -742
rect 2167 -743 2170 -739
rect 2097 -755 2100 -745
rect 2138 -746 2170 -743
rect 2176 -746 2180 -739
rect 2138 -749 2141 -746
rect 2085 -758 2100 -755
rect 2085 -761 2088 -758
rect 2137 -752 2143 -749
rect 2176 -750 2212 -746
rect 2216 -758 2225 -754
rect 2232 -761 2236 -739
rect 2240 -750 2241 -746
rect 2276 -748 2279 -739
rect 2320 -748 2323 -739
rect 2276 -753 2288 -748
rect 2320 -753 2344 -748
rect 2351 -749 2355 -739
rect 2400 -749 2404 -739
rect 2240 -755 2248 -753
rect 2245 -758 2248 -755
rect 2267 -758 2268 -754
rect 2276 -761 2279 -753
rect 2284 -758 2292 -753
rect 2311 -758 2312 -754
rect 2320 -761 2323 -753
rect 2351 -754 2379 -749
rect 2400 -753 2409 -749
rect 2351 -761 2355 -754
rect 2400 -757 2404 -753
rect 2076 -771 2079 -767
rect 2097 -768 2102 -765
rect 2115 -765 2118 -761
rect 2162 -765 2165 -761
rect 2107 -768 2171 -765
rect 2097 -771 2100 -768
rect 2070 -774 2100 -771
rect 2224 -771 2236 -761
rect 2268 -771 2279 -761
rect 2312 -771 2323 -761
rect 2212 -776 2216 -771
rect 2248 -776 2252 -771
rect 2292 -776 2296 -771
rect 2343 -776 2347 -771
rect 2211 -780 2355 -776
rect 2392 -777 2396 -767
rect 2224 -812 2377 -808
rect 2230 -818 2234 -812
rect 2268 -818 2272 -812
rect 2312 -818 2316 -812
rect 2357 -818 2361 -812
rect 2397 -813 2401 -810
rect 2391 -817 2392 -813
rect 2396 -817 2401 -813
rect 2280 -843 2293 -818
rect 2324 -843 2337 -818
rect 2397 -823 2401 -817
rect 2170 -854 2226 -850
rect 2170 -931 2174 -854
rect 2230 -862 2239 -858
rect 2246 -865 2250 -843
rect 2254 -854 2255 -850
rect 2290 -852 2293 -843
rect 2334 -852 2337 -843
rect 2290 -857 2302 -852
rect 2334 -857 2358 -852
rect 2365 -853 2369 -843
rect 2405 -853 2409 -843
rect 2254 -859 2262 -857
rect 2259 -862 2262 -859
rect 2281 -862 2282 -858
rect 2290 -865 2293 -857
rect 2298 -862 2306 -857
rect 2325 -862 2326 -858
rect 2334 -865 2337 -857
rect 2365 -858 2384 -853
rect 2405 -857 2414 -853
rect 2365 -865 2369 -858
rect 2405 -861 2409 -857
rect 2238 -875 2250 -865
rect 2282 -875 2293 -865
rect 2326 -875 2337 -865
rect 2226 -880 2230 -875
rect 2262 -880 2266 -875
rect 2306 -880 2310 -875
rect 2357 -880 2361 -875
rect 2225 -884 2369 -880
rect 2397 -881 2401 -871
rect 2138 -935 2174 -931
rect 2078 -974 2081 -940
rect 2138 -941 2142 -935
rect 2124 -944 2149 -941
rect 2084 -950 2093 -947
rect 2084 -964 2087 -950
rect 2124 -955 2127 -944
rect 2117 -958 2127 -955
rect 2084 -967 2093 -964
rect 2078 -977 2087 -974
rect 2078 -993 2081 -977
rect 2114 -983 2117 -968
rect 2111 -986 2117 -983
rect 2078 -996 2087 -993
rect 2078 -1008 2081 -996
rect 2129 -1005 2132 -965
rect 2140 -976 2143 -954
rect 2146 -970 2149 -944
rect 2168 -946 2171 -940
rect 2377 -941 2530 -937
rect 2164 -949 2171 -946
rect 2152 -970 2155 -968
rect 2146 -973 2155 -970
rect 2152 -974 2155 -973
rect 2140 -979 2148 -976
rect 2074 -1011 2081 -1008
rect 2103 -1008 2132 -1005
rect 2074 -1032 2077 -1011
rect 2103 -1023 2106 -1008
rect 2145 -1011 2148 -979
rect 2168 -993 2171 -949
rect 2383 -947 2387 -941
rect 2421 -947 2425 -941
rect 2465 -947 2469 -941
rect 2510 -947 2514 -941
rect 2558 -942 2562 -939
rect 2552 -946 2553 -942
rect 2557 -946 2562 -942
rect 2433 -972 2446 -947
rect 2477 -972 2490 -947
rect 2558 -952 2562 -946
rect 2307 -983 2379 -979
rect 2164 -996 2171 -993
rect 2168 -1004 2171 -996
rect 2168 -1011 2171 -1009
rect 2145 -1014 2161 -1011
rect 2168 -1014 2177 -1011
rect 2119 -1018 2122 -1017
rect 2119 -1023 2121 -1018
rect 2095 -1026 2109 -1023
rect 2074 -1035 2083 -1032
rect 2074 -1036 2077 -1035
rect 2103 -1044 2106 -1034
rect 2119 -1032 2122 -1023
rect 2115 -1035 2122 -1032
rect 2119 -1041 2122 -1035
rect 2129 -1032 2132 -1017
rect 2158 -1023 2161 -1014
rect 2150 -1026 2164 -1023
rect 2129 -1035 2138 -1032
rect 2129 -1036 2132 -1035
rect 2130 -1041 2132 -1036
rect 2158 -1044 2161 -1034
rect 2174 -1032 2177 -1014
rect 2170 -1035 2177 -1032
rect 2174 -1041 2177 -1035
rect 2247 -1022 2250 -988
rect 2307 -989 2311 -983
rect 2293 -992 2318 -989
rect 2253 -998 2262 -995
rect 2253 -1012 2256 -998
rect 2293 -1003 2296 -992
rect 2286 -1006 2296 -1003
rect 2253 -1015 2262 -1012
rect 2247 -1025 2256 -1022
rect 2247 -1041 2250 -1025
rect 2283 -1031 2286 -1016
rect 2280 -1034 2286 -1031
rect 2247 -1044 2256 -1041
rect 2039 -1253 2043 -1237
rect 2104 -1245 2107 -1049
rect 2158 -1072 2161 -1049
rect 2247 -1056 2250 -1044
rect 2298 -1053 2301 -1013
rect 2309 -1024 2312 -1002
rect 2315 -1018 2318 -992
rect 2337 -994 2340 -988
rect 2383 -991 2392 -987
rect 2399 -994 2403 -972
rect 2407 -983 2408 -979
rect 2443 -981 2446 -972
rect 2487 -981 2490 -972
rect 2443 -986 2455 -981
rect 2487 -986 2511 -981
rect 2518 -982 2522 -972
rect 2566 -982 2570 -972
rect 2407 -988 2415 -986
rect 2412 -991 2415 -988
rect 2434 -991 2435 -987
rect 2443 -994 2446 -986
rect 2451 -991 2459 -986
rect 2478 -991 2479 -987
rect 2487 -994 2490 -986
rect 2518 -987 2545 -982
rect 2566 -986 2575 -982
rect 2518 -994 2522 -987
rect 2566 -990 2570 -986
rect 2333 -997 2340 -994
rect 2321 -1018 2324 -1016
rect 2315 -1021 2324 -1018
rect 2321 -1022 2324 -1021
rect 2309 -1027 2317 -1024
rect 2243 -1059 2250 -1056
rect 2272 -1056 2301 -1053
rect 2157 -1075 2162 -1072
rect 2243 -1080 2246 -1059
rect 2272 -1071 2275 -1056
rect 2314 -1059 2317 -1027
rect 2337 -1041 2340 -997
rect 2391 -1004 2403 -994
rect 2435 -1004 2446 -994
rect 2479 -1004 2490 -994
rect 2379 -1009 2383 -1004
rect 2415 -1009 2419 -1004
rect 2459 -1009 2463 -1004
rect 2510 -1009 2514 -1004
rect 2378 -1013 2522 -1009
rect 2558 -1010 2562 -1000
rect 2333 -1044 2340 -1041
rect 2337 -1052 2340 -1044
rect 2337 -1059 2340 -1057
rect 2314 -1062 2330 -1059
rect 2337 -1062 2346 -1059
rect 2288 -1066 2291 -1065
rect 2288 -1071 2290 -1066
rect 2264 -1074 2278 -1071
rect 2243 -1083 2252 -1080
rect 2243 -1084 2246 -1083
rect 2272 -1092 2275 -1082
rect 2288 -1080 2291 -1071
rect 2284 -1083 2291 -1080
rect 2288 -1089 2291 -1083
rect 2298 -1080 2301 -1065
rect 2327 -1071 2330 -1062
rect 2319 -1074 2333 -1071
rect 2298 -1083 2307 -1080
rect 2298 -1084 2301 -1083
rect 2299 -1089 2301 -1084
rect 2327 -1092 2330 -1082
rect 2343 -1080 2346 -1062
rect 2339 -1083 2346 -1080
rect 2343 -1089 2346 -1083
rect 2096 -1249 2114 -1245
rect 2039 -1257 2056 -1253
rect 2143 -1253 2147 -1237
rect 2134 -1257 2147 -1253
rect 2046 -1258 2050 -1257
rect 2046 -1263 2050 -1262
rect 2007 -1507 2012 -1506
rect 2007 -1512 2012 -1511
rect 1998 -1516 2018 -1512
rect 2007 -1530 2012 -1516
rect 2106 -1520 2110 -1289
rect 2206 -1296 2210 -1276
rect 2273 -1288 2276 -1097
rect 2327 -1102 2330 -1097
rect 2571 -1099 2724 -1095
rect 2577 -1105 2581 -1099
rect 2615 -1105 2619 -1099
rect 2659 -1105 2663 -1099
rect 2704 -1105 2708 -1099
rect 2751 -1100 2755 -1097
rect 2745 -1104 2746 -1100
rect 2750 -1104 2755 -1100
rect 2627 -1130 2640 -1105
rect 2671 -1130 2684 -1105
rect 2751 -1110 2755 -1104
rect 2490 -1141 2573 -1137
rect 2430 -1180 2433 -1146
rect 2490 -1147 2494 -1141
rect 2476 -1150 2501 -1147
rect 2436 -1156 2445 -1153
rect 2436 -1170 2439 -1156
rect 2476 -1161 2479 -1150
rect 2469 -1164 2479 -1161
rect 2436 -1173 2445 -1170
rect 2430 -1183 2439 -1180
rect 2430 -1199 2433 -1183
rect 2466 -1189 2469 -1174
rect 2463 -1192 2469 -1189
rect 2430 -1202 2439 -1199
rect 2430 -1214 2433 -1202
rect 2481 -1211 2484 -1171
rect 2492 -1182 2495 -1160
rect 2498 -1176 2501 -1150
rect 2520 -1152 2523 -1146
rect 2577 -1149 2586 -1145
rect 2593 -1152 2597 -1130
rect 2601 -1141 2602 -1137
rect 2637 -1139 2640 -1130
rect 2681 -1139 2684 -1130
rect 2637 -1144 2649 -1139
rect 2681 -1144 2705 -1139
rect 2712 -1140 2716 -1130
rect 2759 -1140 2763 -1130
rect 2601 -1146 2609 -1144
rect 2606 -1149 2609 -1146
rect 2628 -1149 2629 -1145
rect 2637 -1152 2640 -1144
rect 2645 -1149 2653 -1144
rect 2672 -1149 2673 -1145
rect 2681 -1152 2684 -1144
rect 2712 -1145 2738 -1140
rect 2759 -1144 2768 -1140
rect 2712 -1152 2716 -1145
rect 2759 -1148 2763 -1144
rect 2516 -1155 2523 -1152
rect 2504 -1176 2507 -1174
rect 2498 -1179 2507 -1176
rect 2504 -1180 2507 -1179
rect 2492 -1185 2500 -1182
rect 2426 -1217 2433 -1214
rect 2455 -1214 2484 -1211
rect 2426 -1238 2429 -1217
rect 2455 -1229 2458 -1214
rect 2497 -1217 2500 -1185
rect 2520 -1199 2523 -1155
rect 2585 -1162 2597 -1152
rect 2629 -1162 2640 -1152
rect 2673 -1162 2684 -1152
rect 2573 -1167 2577 -1162
rect 2609 -1167 2613 -1162
rect 2653 -1167 2657 -1162
rect 2704 -1167 2708 -1162
rect 2572 -1171 2716 -1167
rect 2751 -1168 2755 -1158
rect 2516 -1202 2523 -1199
rect 2520 -1210 2523 -1202
rect 2520 -1217 2523 -1215
rect 2497 -1220 2513 -1217
rect 2520 -1220 2529 -1217
rect 2471 -1224 2474 -1223
rect 2471 -1229 2473 -1224
rect 2447 -1232 2461 -1229
rect 2426 -1241 2435 -1238
rect 2426 -1242 2429 -1241
rect 2455 -1250 2458 -1240
rect 2471 -1238 2474 -1229
rect 2467 -1241 2474 -1238
rect 2471 -1247 2474 -1241
rect 2481 -1238 2484 -1223
rect 2510 -1229 2513 -1220
rect 2502 -1232 2516 -1229
rect 2481 -1241 2490 -1238
rect 2481 -1242 2484 -1241
rect 2482 -1247 2484 -1242
rect 2510 -1250 2513 -1240
rect 2526 -1238 2529 -1220
rect 2522 -1241 2529 -1238
rect 2526 -1247 2529 -1241
rect 2263 -1292 2281 -1288
rect 2206 -1300 2223 -1296
rect 2310 -1296 2314 -1276
rect 2301 -1300 2314 -1296
rect 2206 -1307 2210 -1300
rect 2213 -1301 2217 -1300
rect 2213 -1306 2217 -1305
rect 2310 -1307 2314 -1300
rect 2388 -1303 2392 -1287
rect 2456 -1295 2459 -1255
rect 2510 -1258 2513 -1255
rect 2510 -1264 2515 -1258
rect 2445 -1299 2463 -1295
rect 2388 -1307 2405 -1303
rect 2492 -1303 2496 -1287
rect 2483 -1307 2496 -1303
rect 2388 -1315 2392 -1307
rect 2395 -1308 2399 -1307
rect 2395 -1313 2399 -1312
rect 2492 -1315 2496 -1307
rect 2273 -1339 2278 -1333
rect 2181 -1484 2186 -1483
rect 2181 -1489 2186 -1488
rect 2172 -1493 2192 -1489
rect 2181 -1507 2186 -1493
rect 2274 -1497 2278 -1339
rect 2455 -1350 2460 -1346
rect 2456 -1365 2459 -1350
rect 2355 -1480 2360 -1479
rect 2355 -1485 2360 -1484
rect 2346 -1489 2366 -1485
rect 2242 -1501 2278 -1497
rect 2068 -1524 2110 -1520
rect 2106 -1561 2110 -1524
rect 2274 -1551 2278 -1501
rect 2355 -1503 2360 -1489
rect 2455 -1493 2459 -1365
rect 2683 -1378 2704 -1374
rect 2691 -1381 2695 -1378
rect 2685 -1385 2686 -1381
rect 2690 -1385 2695 -1381
rect 2691 -1391 2695 -1385
rect 2732 -1404 2885 -1400
rect 2551 -1445 2556 -1444
rect 2645 -1446 2691 -1441
rect 2699 -1442 2703 -1431
rect 2738 -1410 2742 -1404
rect 2776 -1410 2780 -1404
rect 2820 -1410 2824 -1404
rect 2865 -1410 2869 -1404
rect 2903 -1408 2907 -1405
rect 2788 -1435 2801 -1410
rect 2832 -1435 2845 -1410
rect 2897 -1412 2898 -1408
rect 2902 -1412 2907 -1408
rect 2699 -1446 2734 -1442
rect 2551 -1450 2556 -1449
rect 2542 -1454 2562 -1450
rect 2551 -1468 2556 -1454
rect 2645 -1458 2649 -1446
rect 2699 -1449 2703 -1446
rect 2612 -1462 2649 -1458
rect 2416 -1497 2459 -1493
rect 2455 -1543 2459 -1497
rect 2645 -1535 2649 -1462
rect 2738 -1454 2747 -1450
rect 2754 -1457 2758 -1435
rect 2762 -1446 2763 -1442
rect 2798 -1444 2801 -1435
rect 2842 -1444 2845 -1435
rect 2798 -1449 2810 -1444
rect 2842 -1449 2866 -1444
rect 2873 -1445 2877 -1435
rect 2903 -1418 2907 -1412
rect 2762 -1451 2770 -1449
rect 2767 -1454 2770 -1451
rect 2789 -1454 2790 -1450
rect 2798 -1457 2801 -1449
rect 2806 -1454 2814 -1449
rect 2833 -1454 2834 -1450
rect 2842 -1457 2845 -1449
rect 2873 -1450 2886 -1445
rect 2911 -1448 2915 -1438
rect 2873 -1457 2877 -1450
rect 2911 -1452 2920 -1448
rect 2911 -1456 2915 -1452
rect 2746 -1467 2758 -1457
rect 2790 -1467 2801 -1457
rect 2834 -1467 2845 -1457
rect 2691 -1478 2695 -1469
rect 2734 -1472 2738 -1467
rect 2770 -1472 2774 -1467
rect 2814 -1472 2818 -1467
rect 2865 -1472 2869 -1467
rect 2733 -1476 2877 -1472
rect 2903 -1476 2907 -1466
rect 2683 -1482 2700 -1478
rect 2638 -1539 2649 -1535
rect 2450 -1547 2538 -1543
rect 2273 -1553 2350 -1551
rect 2269 -1555 2350 -1553
rect 2269 -1557 2277 -1555
rect 2101 -1565 2169 -1561
rect 1899 -1783 1918 -1778
rect 1948 -1573 2001 -1569
rect 1948 -1679 1952 -1573
rect 2106 -1675 2110 -1565
rect 2273 -1664 2277 -1557
rect 2454 -1654 2458 -1547
rect 2645 -1644 2649 -1539
rect 2640 -1648 2649 -1644
rect 2448 -1658 2458 -1654
rect 2533 -1656 2540 -1652
rect 2268 -1668 2277 -1664
rect 2342 -1666 2348 -1662
rect 2100 -1679 2110 -1675
rect 2162 -1676 2168 -1672
rect 1994 -1687 2000 -1683
rect 1744 -1799 1767 -1795
rect 1748 -1801 1767 -1799
rect 1744 -1810 1748 -1805
rect 1763 -1810 1767 -1801
rect 1899 -1802 1904 -1783
rect 1915 -1786 1918 -1783
rect 1956 -1781 1960 -1779
rect 1995 -1692 1999 -1687
rect 2162 -1692 2166 -1676
rect 2342 -1692 2346 -1666
rect 2533 -1692 2537 -1656
rect 1995 -1696 2537 -1692
rect 1995 -1781 1999 -1696
rect 2133 -1777 2139 -1773
rect 1956 -1785 2033 -1781
rect 1780 -1806 1804 -1805
rect 1780 -1810 1796 -1806
rect 1800 -1810 1804 -1806
rect 1899 -1807 1939 -1802
rect 1780 -1812 1804 -1810
rect 1786 -1817 1790 -1812
rect 1755 -1838 1759 -1830
rect 1755 -1842 1767 -1838
rect 1763 -1844 1767 -1842
rect 1794 -1844 1798 -1837
rect 1889 -1841 1893 -1825
rect 1934 -1833 1939 -1807
rect 2073 -1812 2077 -1803
rect 2130 -1806 2140 -1804
rect 2145 -1806 2148 -1804
rect 2130 -1808 2148 -1806
rect 2073 -1816 2090 -1812
rect 2177 -1812 2181 -1807
rect 2168 -1816 2181 -1812
rect 2073 -1826 2077 -1816
rect 2080 -1817 2084 -1816
rect 2080 -1822 2084 -1821
rect 2177 -1825 2181 -1816
rect 1924 -1837 1946 -1833
rect 948 -1849 1157 -1845
rect 1162 -1849 1756 -1845
rect 1763 -1848 1787 -1844
rect 1794 -1848 1830 -1844
rect 1889 -1845 1899 -1841
rect 1961 -1841 1965 -1833
rect 948 -1856 1254 -1852
rect 1259 -1856 1745 -1852
rect 1763 -1859 1767 -1848
rect 1794 -1851 1798 -1848
rect 1786 -1865 1790 -1861
rect 1780 -1866 1805 -1865
rect 1780 -1870 1800 -1866
rect 1780 -1871 1805 -1870
rect 1744 -1883 1748 -1879
rect 1744 -1887 1760 -1883
rect 1889 -1886 1893 -1845
rect 1933 -1865 1938 -1844
rect 1956 -1845 1965 -1841
rect 1899 -1868 1956 -1865
rect 1899 -1878 1924 -1868
rect 1939 -1877 1943 -1876
rect 1946 -1876 1956 -1868
rect 1889 -1890 1899 -1886
rect 1745 -1918 1768 -1914
rect 1749 -1920 1768 -1918
rect 1745 -1929 1749 -1924
rect 1764 -1929 1768 -1920
rect 1781 -1925 1805 -1924
rect 1781 -1929 1797 -1925
rect 1801 -1929 1805 -1925
rect 1781 -1931 1805 -1929
rect 1889 -1930 1893 -1890
rect 1961 -1892 1965 -1845
rect 1956 -1896 1965 -1892
rect 1938 -1900 1943 -1896
rect 1933 -1904 1943 -1900
rect 1933 -1909 1938 -1904
rect 1899 -1912 1956 -1909
rect 1899 -1922 1924 -1912
rect 1939 -1921 1943 -1920
rect 1946 -1920 1956 -1912
rect 1787 -1936 1791 -1931
rect 1889 -1934 1899 -1930
rect 1756 -1957 1760 -1949
rect 1756 -1961 1768 -1957
rect 1764 -1963 1768 -1961
rect 1795 -1963 1799 -1956
rect 948 -1968 1460 -1964
rect 1465 -1968 1757 -1964
rect 1764 -1967 1788 -1963
rect 1795 -1967 1842 -1963
rect 948 -1975 1358 -1971
rect 1363 -1975 1746 -1971
rect 1764 -1978 1768 -1967
rect 1795 -1970 1799 -1967
rect 1889 -1968 1893 -1934
rect 1961 -1936 1965 -1896
rect 1956 -1940 1965 -1936
rect 1931 -1948 1935 -1947
rect 1938 -1943 1943 -1940
rect 1938 -1948 1940 -1943
rect 1924 -1956 1956 -1952
rect 1889 -1972 1899 -1968
rect 1939 -1972 1943 -1963
rect 1946 -1964 1956 -1956
rect 1961 -1972 1965 -1940
rect 1889 -1978 1893 -1972
rect 1787 -1984 1791 -1980
rect 1931 -1983 1935 -1976
rect 1956 -1976 1965 -1972
rect 1961 -1977 1965 -1976
rect 1781 -1985 1806 -1984
rect 1781 -1989 1801 -1985
rect 1781 -1990 1806 -1989
rect 1745 -2002 1749 -1998
rect 1745 -2006 1761 -2002
rect 1749 -2026 1772 -2022
rect 1753 -2028 1772 -2026
rect 1749 -2037 1753 -2032
rect 1768 -2037 1772 -2028
rect 1785 -2033 1809 -2032
rect 1785 -2037 1801 -2033
rect 1805 -2037 1809 -2033
rect 1785 -2039 1809 -2037
rect 1791 -2044 1795 -2039
rect 1760 -2065 1764 -2057
rect 1760 -2069 1772 -2065
rect 1768 -2071 1772 -2069
rect 1799 -2071 1803 -2064
rect 948 -2076 1655 -2072
rect 1660 -2076 1761 -2072
rect 1768 -2075 1792 -2071
rect 1799 -2075 1856 -2071
rect 948 -2083 1555 -2079
rect 1562 -2083 1750 -2079
rect 1768 -2086 1772 -2075
rect 1799 -2078 1803 -2075
rect 1791 -2092 1795 -2088
rect 1785 -2093 1810 -2092
rect 1785 -2097 1805 -2093
rect 1785 -2098 1810 -2097
rect 1749 -2110 1753 -2106
rect 1749 -2114 1765 -2110
<< m2contact >>
rect 944 -890 949 -885
rect 942 -919 947 -914
rect 952 -920 957 -915
rect 944 -947 949 -942
rect 944 -991 949 -986
rect 948 -1038 953 -1032
rect 1051 -890 1056 -885
rect 1049 -919 1054 -914
rect 1059 -920 1064 -915
rect 1051 -947 1056 -942
rect 1051 -991 1056 -986
rect 1055 -1038 1060 -1032
rect 1153 -890 1158 -885
rect 1151 -919 1156 -914
rect 1161 -920 1166 -915
rect 1153 -947 1158 -942
rect 1153 -991 1158 -986
rect 1157 -1038 1162 -1032
rect 1250 -890 1255 -885
rect 1248 -919 1253 -914
rect 1258 -920 1263 -915
rect 1250 -947 1255 -942
rect 1250 -991 1255 -986
rect 1254 -1038 1259 -1032
rect 1354 -889 1359 -884
rect 1352 -918 1357 -913
rect 1362 -919 1367 -914
rect 1354 -946 1359 -941
rect 1354 -990 1359 -985
rect 1358 -1037 1363 -1031
rect 1456 -889 1461 -884
rect 1454 -918 1459 -913
rect 1464 -919 1469 -914
rect 1456 -946 1461 -941
rect 1456 -990 1461 -985
rect 1460 -1037 1465 -1031
rect 1552 -889 1557 -884
rect 1550 -918 1555 -913
rect 1560 -919 1565 -914
rect 1552 -946 1557 -941
rect 1552 -990 1557 -985
rect 1556 -1037 1561 -1031
rect 1651 -889 1656 -884
rect 1649 -918 1654 -913
rect 1659 -919 1664 -914
rect 1651 -946 1656 -941
rect 1651 -990 1656 -985
rect 1655 -1036 1660 -1030
rect 1655 -1100 1660 -1095
rect 1697 -1100 1702 -1095
rect 1556 -1153 1561 -1148
rect 1697 -1154 1702 -1149
rect 1811 -1174 1816 -1169
rect 1460 -1231 1465 -1226
rect 1698 -1232 1703 -1227
rect 1358 -1285 1363 -1280
rect 1698 -1286 1703 -1281
rect 1811 -1304 1816 -1299
rect 1254 -1375 1259 -1370
rect 1701 -1376 1706 -1371
rect 1157 -1429 1162 -1424
rect 1701 -1430 1706 -1425
rect 1815 -1450 1820 -1445
rect 1055 -1501 1060 -1496
rect 1708 -1501 1713 -1496
rect 948 -1555 953 -1550
rect 1708 -1555 1713 -1550
rect 1822 -1577 1827 -1572
rect 1055 -1740 1060 -1735
rect 948 -1748 953 -1743
rect 1817 -1740 1822 -1735
rect 2062 -705 2067 -700
rect 1989 -758 1994 -753
rect 2062 -759 2067 -754
rect 2211 -758 2216 -753
rect 2241 -750 2246 -745
rect 2240 -760 2245 -755
rect 2268 -758 2273 -753
rect 2312 -758 2317 -753
rect 2379 -754 2386 -749
rect 2225 -862 2230 -857
rect 2255 -854 2260 -849
rect 2254 -864 2259 -859
rect 2282 -862 2287 -857
rect 2326 -862 2331 -857
rect 2384 -858 2391 -853
rect 2103 -1049 2108 -1044
rect 2157 -1049 2162 -1044
rect 2378 -991 2383 -986
rect 2408 -983 2413 -978
rect 2407 -993 2412 -988
rect 2435 -991 2440 -986
rect 2479 -991 2484 -986
rect 2545 -987 2551 -982
rect 2157 -1080 2162 -1075
rect 2272 -1097 2277 -1092
rect 2326 -1097 2331 -1092
rect 2106 -1289 2111 -1283
rect 2327 -1108 2333 -1102
rect 2572 -1149 2577 -1144
rect 2602 -1141 2607 -1136
rect 2601 -1151 2606 -1146
rect 2629 -1149 2634 -1144
rect 2673 -1149 2678 -1144
rect 2738 -1145 2745 -1140
rect 2455 -1255 2460 -1250
rect 2509 -1255 2514 -1250
rect 2510 -1270 2515 -1264
rect 2273 -1333 2278 -1325
rect 2455 -1346 2460 -1340
rect 2733 -1454 2738 -1449
rect 2763 -1446 2768 -1441
rect 2762 -1456 2767 -1451
rect 2790 -1454 2795 -1449
rect 2834 -1454 2839 -1449
rect 1915 -1791 1920 -1786
rect 2140 -1806 2145 -1801
rect 1157 -1849 1162 -1844
rect 1830 -1848 1835 -1843
rect 1254 -1857 1259 -1852
rect 1938 -1876 1943 -1871
rect 1938 -1920 1943 -1915
rect 1460 -1968 1465 -1963
rect 1842 -1967 1848 -1961
rect 1358 -1976 1363 -1971
rect 1930 -1947 1935 -1942
rect 1940 -1948 1945 -1943
rect 1938 -1977 1943 -1972
rect 1655 -2076 1660 -2071
rect 1856 -2075 1861 -2069
rect 1555 -2084 1562 -2079
<< pm12contact >>
rect 1753 -1117 1758 -1112
rect 1762 -1118 1767 -1113
rect 1754 -1249 1759 -1244
rect 1763 -1250 1768 -1245
rect 1757 -1393 1762 -1388
rect 1766 -1394 1771 -1389
rect 1764 -1518 1769 -1513
rect 1773 -1519 1778 -1514
rect 2118 -722 2123 -717
rect 2127 -723 2132 -718
rect 2392 -754 2397 -749
rect 2397 -858 2402 -853
rect 2121 -984 2126 -979
rect 2120 -993 2125 -988
rect 2290 -1032 2295 -1027
rect 2289 -1041 2294 -1036
rect 2558 -987 2563 -982
rect 2106 -1257 2111 -1252
rect 2085 -1517 2091 -1511
rect 2473 -1190 2478 -1185
rect 2472 -1199 2477 -1194
rect 2751 -1145 2756 -1140
rect 2273 -1300 2278 -1295
rect 2455 -1307 2460 -1302
rect 2259 -1494 2265 -1488
rect 2433 -1490 2439 -1484
rect 2629 -1455 2635 -1449
rect 2903 -1453 2908 -1448
rect 2526 -1540 2531 -1535
rect 2338 -1548 2343 -1543
rect 2157 -1558 2162 -1553
rect 1989 -1566 1994 -1561
rect 2528 -1649 2533 -1644
rect 2336 -1659 2341 -1654
rect 2156 -1669 2161 -1664
rect 1988 -1680 1993 -1675
rect 2140 -1785 2145 -1780
rect 1948 -1791 1953 -1786
rect 2140 -1816 2145 -1811
<< metal2 >>
rect 2241 -700 2272 -697
rect 2063 -711 2066 -705
rect 2063 -714 2100 -711
rect 2097 -717 2100 -714
rect 2097 -720 2118 -717
rect 2127 -733 2130 -723
rect 2064 -736 2130 -733
rect 2064 -754 2067 -736
rect 2241 -745 2245 -700
rect 2268 -753 2272 -700
rect 944 -876 948 -864
rect 1051 -876 1055 -864
rect 1153 -876 1157 -864
rect 1250 -876 1254 -864
rect 1354 -875 1358 -863
rect 1456 -875 1460 -863
rect 1552 -875 1556 -863
rect 1651 -875 1655 -863
rect 917 -882 948 -876
rect 917 -915 920 -882
rect 944 -885 948 -882
rect 1024 -882 1055 -876
rect 917 -919 942 -915
rect 1024 -915 1027 -882
rect 1051 -885 1055 -882
rect 1126 -882 1157 -876
rect 917 -986 920 -919
rect 957 -919 1005 -915
rect 1002 -942 1005 -919
rect 949 -946 1005 -942
rect 1024 -919 1049 -915
rect 1126 -915 1129 -882
rect 1153 -885 1157 -882
rect 1223 -882 1254 -876
rect 1024 -986 1027 -919
rect 1064 -919 1112 -915
rect 1109 -942 1112 -919
rect 1056 -946 1112 -942
rect 1126 -919 1151 -915
rect 1223 -915 1226 -882
rect 1250 -885 1254 -882
rect 1327 -881 1358 -875
rect 1327 -914 1330 -881
rect 1354 -884 1358 -881
rect 1429 -881 1460 -875
rect 1126 -986 1129 -919
rect 1166 -919 1214 -915
rect 1211 -942 1214 -919
rect 1158 -946 1214 -942
rect 1223 -919 1248 -915
rect 1223 -986 1226 -919
rect 1263 -919 1311 -915
rect 1308 -942 1311 -919
rect 1255 -946 1311 -942
rect 1327 -918 1352 -914
rect 1429 -914 1432 -881
rect 1456 -884 1460 -881
rect 1525 -881 1556 -875
rect 1327 -985 1330 -918
rect 1367 -918 1415 -914
rect 1412 -941 1415 -918
rect 1359 -945 1415 -941
rect 1429 -918 1454 -914
rect 1525 -914 1528 -881
rect 1552 -884 1556 -881
rect 1624 -881 1655 -875
rect 1429 -985 1432 -918
rect 1469 -918 1517 -914
rect 1514 -941 1517 -918
rect 1461 -945 1517 -941
rect 1525 -918 1550 -914
rect 1624 -914 1627 -881
rect 1651 -884 1655 -881
rect 1525 -985 1528 -918
rect 1565 -918 1613 -914
rect 1610 -941 1613 -918
rect 1557 -945 1613 -941
rect 1624 -918 1649 -914
rect 1624 -985 1627 -918
rect 1664 -918 1712 -914
rect 1709 -941 1712 -918
rect 1656 -945 1712 -941
rect 917 -991 944 -986
rect 1024 -991 1051 -986
rect 1126 -991 1153 -986
rect 1223 -991 1250 -986
rect 1327 -990 1354 -985
rect 1429 -990 1456 -985
rect 1525 -990 1552 -985
rect 1624 -990 1651 -985
rect 917 -995 920 -991
rect 1024 -995 1027 -991
rect 1126 -995 1129 -991
rect 1223 -995 1226 -991
rect 1327 -994 1330 -990
rect 1429 -994 1432 -990
rect 1525 -994 1528 -990
rect 1624 -994 1627 -990
rect 1055 -1032 1060 -1031
rect 1254 -1032 1259 -1029
rect 948 -1550 953 -1038
rect 948 -1743 953 -1555
rect 948 -2083 953 -1748
rect 1055 -1496 1060 -1038
rect 1055 -1735 1060 -1501
rect 1055 -2083 1060 -1740
rect 1157 -1424 1162 -1038
rect 1157 -1844 1162 -1429
rect 1157 -2083 1162 -1849
rect 1254 -1370 1259 -1038
rect 1254 -1852 1259 -1375
rect 1254 -2083 1259 -1857
rect 1358 -1031 1363 -1028
rect 1358 -1280 1363 -1037
rect 1358 -1971 1363 -1285
rect 1358 -2083 1363 -1976
rect 1460 -1031 1465 -1028
rect 1460 -1226 1465 -1037
rect 1460 -1963 1465 -1231
rect 1460 -2083 1465 -1968
rect 1556 -1031 1561 -1028
rect 1556 -1148 1561 -1037
rect 1556 -2079 1561 -1153
rect 1655 -1030 1660 -1028
rect 1655 -1095 1660 -1036
rect 1655 -2071 1660 -1100
rect 1698 -1106 1701 -1100
rect 1698 -1109 1735 -1106
rect 1732 -1112 1735 -1109
rect 1732 -1115 1753 -1112
rect 1762 -1128 1765 -1118
rect 1699 -1131 1765 -1128
rect 1699 -1149 1702 -1131
rect 1816 -1174 1871 -1169
rect 1699 -1238 1702 -1232
rect 1699 -1241 1736 -1238
rect 1733 -1244 1736 -1241
rect 1733 -1247 1754 -1244
rect 1763 -1260 1766 -1250
rect 1700 -1263 1766 -1260
rect 1700 -1281 1703 -1263
rect 1816 -1304 1859 -1299
rect 1702 -1382 1705 -1376
rect 1702 -1385 1739 -1382
rect 1736 -1388 1739 -1385
rect 1736 -1391 1757 -1388
rect 1766 -1404 1769 -1394
rect 1703 -1407 1769 -1404
rect 1703 -1425 1706 -1407
rect 1820 -1449 1838 -1445
rect 1709 -1507 1712 -1501
rect 1709 -1510 1746 -1507
rect 1743 -1513 1746 -1510
rect 1743 -1516 1764 -1513
rect 1773 -1529 1776 -1519
rect 1710 -1532 1776 -1529
rect 1710 -1550 1713 -1532
rect 1822 -1613 1827 -1577
rect 1834 -1603 1838 -1449
rect 1854 -1593 1859 -1304
rect 1866 -1578 1871 -1174
rect 1989 -1553 1994 -758
rect 2190 -758 2211 -754
rect 2202 -782 2208 -758
rect 2386 -754 2392 -749
rect 2241 -782 2245 -760
rect 2312 -782 2317 -758
rect 2202 -785 2321 -782
rect 2255 -804 2286 -801
rect 2255 -849 2259 -804
rect 2282 -857 2286 -804
rect 2204 -862 2225 -858
rect 2216 -886 2222 -862
rect 2391 -858 2397 -853
rect 2255 -886 2259 -864
rect 2326 -886 2331 -862
rect 2216 -889 2335 -886
rect 2408 -933 2439 -930
rect 2408 -978 2412 -933
rect 2126 -984 2139 -981
rect 2120 -1011 2123 -993
rect 2114 -1014 2123 -1011
rect 2114 -1045 2117 -1014
rect 2108 -1048 2117 -1045
rect 2136 -1044 2139 -984
rect 2435 -986 2439 -933
rect 2357 -991 2378 -987
rect 2369 -1015 2375 -991
rect 2551 -987 2558 -982
rect 2408 -1015 2412 -993
rect 2479 -1015 2484 -991
rect 2369 -1018 2488 -1015
rect 2295 -1032 2308 -1029
rect 2136 -1047 2157 -1044
rect 2289 -1059 2292 -1041
rect 2283 -1062 2292 -1059
rect 2106 -1283 2111 -1257
rect 2085 -1511 2091 -1507
rect 2157 -1543 2162 -1080
rect 2283 -1093 2286 -1062
rect 2277 -1096 2286 -1093
rect 2305 -1092 2308 -1032
rect 2602 -1091 2633 -1088
rect 2305 -1095 2326 -1092
rect 2333 -1108 2342 -1104
rect 2273 -1325 2278 -1300
rect 2259 -1488 2265 -1484
rect 2338 -1534 2342 -1108
rect 2602 -1136 2606 -1091
rect 2629 -1144 2633 -1091
rect 2551 -1149 2572 -1145
rect 2563 -1173 2569 -1149
rect 2745 -1145 2751 -1140
rect 2602 -1173 2606 -1151
rect 2673 -1173 2678 -1149
rect 2563 -1176 2682 -1173
rect 2478 -1190 2491 -1187
rect 2472 -1217 2475 -1199
rect 2466 -1220 2475 -1217
rect 2466 -1251 2469 -1220
rect 2460 -1254 2469 -1251
rect 2488 -1250 2491 -1190
rect 2488 -1253 2509 -1250
rect 2455 -1340 2460 -1307
rect 2510 -1359 2515 -1270
rect 2510 -1364 2531 -1359
rect 2510 -1365 2515 -1364
rect 2433 -1484 2439 -1480
rect 2526 -1522 2531 -1364
rect 2763 -1396 2794 -1393
rect 2629 -1449 2635 -1445
rect 2763 -1441 2767 -1396
rect 2790 -1449 2794 -1396
rect 2712 -1454 2733 -1450
rect 2724 -1478 2730 -1454
rect 2894 -1453 2903 -1448
rect 2763 -1478 2767 -1456
rect 2834 -1478 2839 -1454
rect 2724 -1481 2843 -1478
rect 1979 -1558 1994 -1553
rect 1979 -1578 1984 -1558
rect 1989 -1561 1994 -1558
rect 2148 -1548 2162 -1543
rect 1866 -1583 1984 -1578
rect 2148 -1593 2153 -1548
rect 2157 -1553 2162 -1548
rect 2329 -1538 2342 -1534
rect 1854 -1598 2153 -1593
rect 2329 -1603 2333 -1538
rect 2338 -1539 2342 -1538
rect 2513 -1527 2531 -1522
rect 2338 -1543 2343 -1539
rect 1834 -1607 2333 -1603
rect 2513 -1613 2518 -1527
rect 2526 -1535 2531 -1527
rect 1822 -1618 2518 -1613
rect 1817 -1642 2533 -1637
rect 1817 -1735 1822 -1642
rect 2528 -1644 2533 -1642
rect 1830 -1652 2341 -1647
rect 1830 -1843 1835 -1652
rect 2336 -1654 2341 -1652
rect 1842 -1663 2161 -1657
rect 1842 -1961 1848 -1663
rect 2156 -1664 2161 -1663
rect 1856 -1672 1993 -1667
rect 1856 -2069 1861 -1672
rect 1988 -1675 1993 -1672
rect 1920 -1791 1948 -1786
rect 2140 -1791 2145 -1785
rect 2140 -1801 2145 -1796
rect 2140 -1819 2145 -1816
rect 1967 -1871 1970 -1867
rect 1943 -1876 1970 -1871
rect 1882 -1920 1938 -1916
rect 1882 -1943 1886 -1920
rect 1882 -1947 1930 -1943
rect 1967 -1943 1970 -1876
rect 1945 -1947 1970 -1943
rect 1939 -1980 1943 -1977
rect 1967 -1980 1970 -1947
rect 1939 -1986 1970 -1980
rect 1939 -1998 1943 -1986
rect 1655 -2083 1660 -2076
<< m3contact >>
rect 2085 -1507 2091 -1501
rect 2259 -1484 2265 -1478
rect 2433 -1480 2439 -1474
rect 2629 -1445 2635 -1439
rect 2140 -1796 2145 -1791
<< m123contact >>
rect 2070 -674 2075 -669
rect 2070 -727 2075 -722
rect 2088 -723 2093 -718
rect 1705 -1069 1710 -1064
rect 1705 -1122 1710 -1117
rect 1723 -1118 1728 -1113
rect 1737 -1163 1742 -1158
rect 1706 -1201 1711 -1196
rect 1706 -1254 1711 -1249
rect 1724 -1250 1729 -1245
rect 1738 -1295 1743 -1290
rect 1709 -1345 1714 -1340
rect 1709 -1398 1714 -1393
rect 1727 -1394 1732 -1389
rect 1741 -1439 1746 -1434
rect 1716 -1470 1721 -1465
rect 1716 -1523 1721 -1518
rect 1734 -1519 1739 -1514
rect 1748 -1564 1753 -1559
rect 2102 -768 2107 -763
rect 2072 -1041 2077 -1036
rect 2121 -1023 2126 -1018
rect 2125 -1041 2130 -1036
rect 2166 -1009 2171 -1004
rect 2241 -1089 2246 -1084
rect 2290 -1071 2295 -1066
rect 2294 -1089 2299 -1084
rect 2335 -1057 2340 -1052
rect 2424 -1247 2429 -1242
rect 2473 -1229 2478 -1224
rect 2477 -1247 2482 -1242
rect 2518 -1215 2523 -1210
<< metal3 >>
rect 2070 -722 2073 -674
rect 2093 -723 2105 -720
rect 2102 -763 2105 -723
rect 2123 -1009 2166 -1006
rect 2123 -1018 2126 -1009
rect 2077 -1041 2125 -1038
rect 2292 -1057 2335 -1054
rect 2292 -1066 2295 -1057
rect 1705 -1117 1708 -1069
rect 2246 -1089 2294 -1086
rect 1728 -1118 1740 -1115
rect 1737 -1158 1740 -1118
rect 1706 -1249 1709 -1201
rect 2475 -1215 2518 -1212
rect 2475 -1224 2478 -1215
rect 2429 -1247 2477 -1244
rect 1729 -1250 1741 -1247
rect 1738 -1290 1741 -1250
rect 1709 -1393 1712 -1345
rect 1732 -1394 1744 -1391
rect 1741 -1434 1744 -1394
rect 2085 -1414 2635 -1409
rect 1716 -1518 1719 -1470
rect 2085 -1501 2091 -1414
rect 2259 -1478 2265 -1414
rect 1739 -1519 1751 -1516
rect 1748 -1559 1751 -1519
rect 2297 -1791 2302 -1414
rect 2433 -1474 2439 -1414
rect 2629 -1439 2635 -1414
rect 2145 -1796 2302 -1791
<< labels >>
rlabel metal1 2103 -1679 2108 -1675 3 pdr1
rlabel metal2 1988 -1675 1993 -1671 3 gen_1
rlabel metal1 1948 -1676 1952 -1671 1 prop1_car0
rlabel metal2 1944 -1791 1948 -1786 1 carry_0
rlabel metal1 1956 -1785 1960 -1780 1 clock_car0
rlabel metal1 2025 -1785 2030 -1781 7 clock_car0
rlabel metal2 2140 -1789 2145 -1785 7 clock_in
rlabel metal1 2134 -1777 2139 -1773 7 gnd!
rlabel metal1 1994 -1687 1999 -1683 3 clock_car0
rlabel metal1 2105 -1565 2109 -1561 3 pdr1
rlabel metal2 1989 -1561 1994 -1557 4 prop_1
rlabel metal1 1995 -1573 2000 -1569 3 prop1_car0
rlabel metal1 1998 -1516 2003 -1512 3 vdd!
rlabel m3contact 2085 -1507 2091 -1501 6 clock_in
rlabel metal1 2077 -1524 2082 -1520 7 pdr1
rlabel metal1 2162 -1676 2167 -1672 3 clock_car0
rlabel metal2 2156 -1664 2161 -1660 3 gen_2
rlabel metal1 2271 -1668 2276 -1664 3 pdr2
rlabel metal1 2272 -1557 2277 -1553 3 pdr2
rlabel metal2 2157 -1553 2162 -1549 3 prop_2
rlabel metal1 2163 -1565 2168 -1561 3 pdr1
rlabel metal1 2172 -1493 2177 -1489 3 vdd!
rlabel m3contact 2259 -1484 2265 -1478 7 clock_in
rlabel metal1 2252 -1501 2256 -1497 7 pdr2
rlabel metal1 2342 -1666 2347 -1662 3 clock_car0
rlabel metal2 2336 -1654 2341 -1650 3 gen_3
rlabel metal1 2451 -1658 2456 -1654 3 pdr3
rlabel metal1 2643 -1648 2648 -1644 3 pdr4
rlabel metal2 2528 -1644 2533 -1640 3 gen_4
rlabel metal1 2534 -1656 2539 -1652 1 clock_car0
rlabel metal1 2453 -1547 2458 -1543 3 pdr3
rlabel metal2 2338 -1543 2343 -1539 3 prop_3
rlabel metal1 2344 -1555 2349 -1551 3 pdr2
rlabel metal1 2641 -1539 2646 -1535 3 pdr4
rlabel metal2 2526 -1535 2531 -1531 3 prop_4
rlabel metal1 2532 -1547 2537 -1543 3 pdr3
rlabel metal1 2346 -1489 2351 -1485 3 vdd!
rlabel m3contact 2433 -1480 2439 -1474 7 clock_in
rlabel metal1 2426 -1497 2430 -1493 7 pdr3
rlabel metal1 2542 -1454 2547 -1450 3 vdd!
rlabel m3contact 2629 -1444 2635 -1439 7 clock_in
rlabel metal1 2622 -1462 2626 -1458 7 pdr4
rlabel metal1 2699 -1446 2703 -1441 1 c4
rlabel metal1 2692 -1378 2697 -1374 5 vdd!
rlabel metal1 2696 -1482 2700 -1478 1 gnd!
rlabel metal1 2742 -1474 2745 -1473 1 gnd
rlabel metal1 2748 -1402 2750 -1401 5 vdd
rlabel metal2 2729 -1453 2729 -1453 1 clk_org
rlabel metal1 2729 -1444 2729 -1444 1 c4
rlabel metal1 2884 -1447 2884 -1447 7 q_c4
rlabel metal1 2906 -1409 2906 -1409 5 vdd!
rlabel metal1 2906 -1473 2906 -1473 1 gnd!
rlabel metal2 2896 -1450 2896 -1450 1 q_c4
rlabel metal1 2918 -1451 2918 -1451 7 iq_c4
rlabel metal1 2177 -1811 2181 -1807 7 gnd!
rlabel metal1 2073 -1815 2077 -1810 3 vdd!
rlabel metal2 2140 -1819 2145 -1816 7 clk_org
rlabel metal1 2140 -1808 2145 -1804 7 clock_in
rlabel metal1 2408 -751 2408 -751 1 iq_s1
rlabel m2contact 2385 -752 2385 -752 1 q_s1
rlabel metal1 2395 -774 2395 -774 1 gnd!
rlabel metal1 2395 -710 2395 -710 5 vdd!
rlabel metal1 2362 -751 2362 -751 7 q_s1
rlabel metal1 2207 -748 2207 -748 1 s1
rlabel metal2 2207 -757 2207 -757 1 clk_org
rlabel metal1 2226 -706 2228 -705 5 vdd
rlabel metal1 2220 -778 2223 -777 1 gnd
rlabel metal1 2179 -737 2179 -737 1 s1
rlabel metal1 2060 -756 2060 -756 1 prop_1
rlabel metal1 2060 -702 2060 -702 1 carry_0
rlabel metal1 2083 -728 2086 -726 1 vdd
rlabel metal1 2082 -674 2085 -672 5 vdd
rlabel metal1 2086 -718 2087 -716 1 gnd
rlabel metal1 2138 -768 2141 -766 1 gnd
rlabel metal1 2088 -774 2092 -771 1 gnd
rlabel metal1 1759 -2025 1759 -2025 5 vdd
rlabel metal1 1760 -2112 1760 -2112 1 gnd
rlabel metal1 1792 -2094 1792 -2094 1 gnd
rlabel metal1 1789 -2037 1789 -2037 5 vdd
rlabel metal1 1744 -2074 1744 -2074 3 q_a1
rlabel metal1 1746 -2081 1746 -2081 3 q_b1
rlabel metal1 1808 -2074 1808 -2074 1 gen_1
rlabel metal1 1755 -1917 1755 -1917 5 vdd
rlabel metal1 1756 -2004 1756 -2004 1 gnd
rlabel metal1 1788 -1986 1788 -1986 1 gnd
rlabel metal1 1785 -1929 1785 -1929 5 vdd
rlabel metal1 1741 -1967 1741 -1967 1 q_a2
rlabel metal1 1741 -1974 1741 -1974 1 q_b2
rlabel metal1 1804 -1965 1804 -1965 1 gen_2
rlabel metal1 1754 -1798 1754 -1798 5 vdd
rlabel metal1 1755 -1885 1755 -1885 1 gnd
rlabel metal1 1787 -1867 1787 -1867 1 gnd
rlabel metal1 1784 -1810 1784 -1810 5 vdd
rlabel metal1 1739 -1848 1739 -1848 1 q_b3
rlabel metal1 1741 -1855 1741 -1855 1 q_a3
rlabel metal1 1802 -1846 1802 -1846 1 gen_3
rlabel metal1 1754 -1689 1754 -1689 5 vdd
rlabel metal1 1755 -1776 1755 -1776 1 gnd
rlabel metal1 1787 -1758 1787 -1758 1 gnd
rlabel metal1 1784 -1701 1784 -1701 5 vdd
rlabel metal1 1739 -1738 1739 -1738 3 q_a4
rlabel metal1 1739 -1744 1739 -1744 3 q_b4
rlabel metal1 1802 -1737 1802 -1737 1 gen_4
rlabel metal1 1814 -1263 1814 -1263 1 prop_2
rlabel metal1 1696 -1284 1696 -1284 3 q_b2
rlabel metal1 1696 -1229 1696 -1229 3 q_a2
rlabel metal1 1719 -1255 1722 -1253 1 vdd
rlabel metal1 1718 -1201 1721 -1199 5 vdd
rlabel metal1 1722 -1245 1723 -1243 1 gnd
rlabel metal1 1774 -1295 1777 -1293 1 gnd
rlabel metal1 1724 -1301 1728 -1298 1 gnd
rlabel metal1 1727 -1445 1731 -1442 1 gnd
rlabel metal1 1777 -1439 1780 -1437 1 gnd
rlabel metal1 1725 -1389 1726 -1387 1 gnd
rlabel metal1 1721 -1345 1724 -1343 5 vdd
rlabel metal1 1722 -1399 1725 -1397 1 vdd
rlabel metal1 1700 -1373 1700 -1373 1 q_a3
rlabel metal1 1700 -1427 1700 -1427 1 q_b3
rlabel metal1 1817 -1408 1817 -1408 1 prop_3
rlabel metal1 1734 -1570 1738 -1567 1 gnd
rlabel metal1 1784 -1564 1787 -1562 1 gnd
rlabel metal1 1732 -1514 1733 -1512 1 gnd
rlabel metal1 1728 -1470 1731 -1468 5 vdd
rlabel metal1 1729 -1524 1732 -1522 1 vdd
rlabel metal1 1706 -1499 1706 -1499 1 q_a4
rlabel metal1 1706 -1552 1706 -1552 1 q_b4
rlabel metal1 1825 -1533 1825 -1533 1 prop_4
rlabel metal1 1811 -1132 1811 -1132 1 prop_1
rlabel metal1 1695 -1151 1695 -1151 1 q_b1
rlabel metal1 1695 -1097 1695 -1097 1 q_a1
rlabel metal1 1718 -1123 1721 -1121 1 vdd
rlabel metal1 1717 -1069 1720 -1067 5 vdd
rlabel metal1 1721 -1113 1722 -1111 1 gnd
rlabel metal1 1773 -1163 1776 -1161 1 gnd
rlabel metal1 1723 -1169 1727 -1166 1 gnd
rlabel metal1 1962 -1968 1963 -1965 7 gnd
rlabel metal1 1890 -1962 1891 -1960 3 vdd
rlabel metal2 1942 -1981 1942 -1981 7 clk_org
rlabel metal1 1933 -1982 1933 -1982 7 cin
rlabel metal1 1937 -1825 1937 -1825 7 carry_0
rlabel metal1 1562 -880 1562 -880 3 b1
rlabel metal2 1553 -880 1553 -880 3 clk_org
rlabel metal1 1604 -901 1605 -899 7 vdd
rlabel metal1 1532 -896 1533 -893 3 gnd
rlabel m2contact 1658 -1035 1658 -1035 3 q_a1
rlabel metal1 1661 -880 1661 -880 3 a1
rlabel metal2 1652 -880 1652 -880 3 clk_org
rlabel metal1 1703 -901 1704 -899 7 vdd
rlabel metal1 1631 -896 1632 -893 3 gnd
rlabel m2contact 1462 -1035 1462 -1035 3 q_a2
rlabel metal1 1466 -880 1466 -880 3 a2
rlabel metal2 1457 -880 1457 -880 3 clk_org
rlabel metal1 1508 -901 1509 -899 7 vdd
rlabel metal1 1436 -896 1437 -893 3 gnd
rlabel m2contact 1360 -1034 1360 -1034 3 q_b2
rlabel metal1 1364 -881 1364 -881 3 b2
rlabel metal2 1355 -880 1355 -880 3 clk_org
rlabel metal1 1406 -901 1407 -899 7 vdd
rlabel metal1 1334 -896 1335 -893 3 gnd
rlabel m2contact 1256 -1035 1256 -1035 3 q_a3
rlabel metal1 1260 -881 1260 -881 3 a3
rlabel metal2 1251 -881 1251 -881 3 clk_org
rlabel metal1 1302 -902 1303 -900 7 vdd
rlabel metal1 1230 -897 1231 -894 3 gnd
rlabel m2contact 1160 -1037 1160 -1037 3 q_b3
rlabel metal1 1163 -882 1163 -882 3 b3
rlabel metal2 1154 -881 1154 -881 3 clk_org
rlabel metal1 1205 -902 1206 -900 7 vdd
rlabel metal1 1133 -897 1134 -894 3 gnd
rlabel m2contact 1057 -1036 1057 -1036 3 q_a4
rlabel metal1 1062 -881 1062 -881 3 a4
rlabel metal2 1052 -881 1052 -881 3 clk_org
rlabel metal1 1103 -902 1104 -900 7 vdd
rlabel metal1 1031 -897 1032 -894 3 gnd
rlabel m2contact 951 -1036 951 -1036 3 q_b4
rlabel metal1 954 -881 954 -881 3 b4
rlabel metal2 945 -881 945 -881 3 clk_org
rlabel metal1 996 -902 997 -900 7 vdd
rlabel metal1 924 -897 925 -894 3 gnd
rlabel m2contact 1559 -1035 1559 -1035 3 q_b1
rlabel metal1 2458 -1257 2458 -1257 7 c3
rlabel metal1 2511 -1257 2511 -1257 7 prop_4
rlabel metal1 2492 -1139 2492 -1139 7 s4
rlabel metal1 2481 -1234 2483 -1231 7 vdd
rlabel metal1 2427 -1235 2429 -1232 3 vdd
rlabel metal1 2471 -1231 2473 -1230 7 gnd
rlabel metal1 2521 -1179 2523 -1176 7 gnd
rlabel metal1 2526 -1229 2529 -1225 7 gnd
rlabel metal1 2581 -1169 2584 -1168 1 gnd
rlabel metal1 2587 -1097 2589 -1096 5 vdd
rlabel metal2 2568 -1148 2568 -1148 1 clk_org
rlabel metal1 2568 -1139 2568 -1139 1 s4
rlabel metal1 2722 -1143 2722 -1143 1 q_s4
rlabel metal1 2754 -1101 2754 -1101 5 vdd!
rlabel metal1 2754 -1165 2754 -1165 1 gnd!
rlabel metal2 2745 -1142 2745 -1142 1 q_s4
rlabel metal1 2766 -1142 2766 -1142 1 iq_s4
rlabel metal2 2455 -1310 2460 -1307 7 pdr3
rlabel metal1 2455 -1299 2460 -1295 7 c3
rlabel metal1 2388 -1307 2392 -1303 3 vdd!
rlabel metal1 2492 -1303 2496 -1299 7 gnd!
rlabel metal1 2174 -1023 2177 -1019 7 gnd
rlabel metal1 2169 -973 2171 -970 7 gnd
rlabel metal1 2119 -1025 2121 -1024 7 gnd
rlabel metal1 2075 -1029 2077 -1026 3 vdd
rlabel metal1 2129 -1028 2131 -1025 7 vdd
rlabel metal1 2106 -1050 2106 -1050 7 c1
rlabel metal1 2160 -1051 2160 -1051 7 prop_2
rlabel metal1 2141 -932 2141 -932 5 s2
rlabel metal1 2234 -882 2237 -881 1 gnd
rlabel metal1 2240 -810 2242 -809 5 vdd
rlabel metal2 2221 -861 2221 -861 1 clk_org
rlabel metal1 2222 -852 2222 -852 1 s2
rlabel metal1 2375 -856 2375 -856 1 q_s2
rlabel metal1 2400 -814 2400 -814 5 vdd!
rlabel metal1 2400 -878 2400 -878 1 gnd!
rlabel metal2 2391 -856 2391 -856 1 q_s2
rlabel metal1 2412 -855 2412 -855 1 iq_s2
rlabel metal1 2343 -1071 2346 -1067 7 gnd
rlabel metal1 2338 -1021 2340 -1018 7 gnd
rlabel metal1 2288 -1073 2290 -1072 7 gnd
rlabel metal1 2244 -1077 2246 -1074 3 vdd
rlabel metal1 2298 -1076 2300 -1073 7 vdd
rlabel metal1 2274 -1099 2274 -1099 7 c2
rlabel metal1 2309 -980 2309 -980 7 s3
rlabel metal1 2329 -1101 2329 -1101 7 prop_3
rlabel metal1 2387 -1011 2390 -1010 1 gnd
rlabel metal1 2393 -939 2395 -938 5 vdd
rlabel metal2 2374 -990 2374 -990 1 clk_org
rlabel metal1 2374 -981 2374 -981 1 s3
rlabel metal1 2529 -984 2529 -984 1 q_s3
rlabel metal1 2561 -943 2561 -943 5 vdd!
rlabel metal1 2561 -1007 2561 -1007 1 gnd!
rlabel metal2 2551 -985 2551 -985 1 q_s3
rlabel metal1 2573 -984 2573 -984 1 iq_s3
rlabel metal1 2143 -1248 2147 -1244 7 gnd!
rlabel metal1 2039 -1257 2043 -1253 3 vdd!
rlabel metal1 2106 -1249 2111 -1245 7 c1
rlabel metal2 2106 -1260 2111 -1257 7 pdr1
rlabel metal1 2310 -1289 2314 -1285 7 gnd!
rlabel metal1 2206 -1300 2210 -1296 3 vdd!
rlabel metal1 2273 -1292 2278 -1288 7 c2
rlabel metal2 2273 -1303 2278 -1300 7 pdr2
<< end >>
